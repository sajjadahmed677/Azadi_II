magic
tech sky130A
magscale 1 2
<<<<<<< HEAD
timestamp 1640101730
=======
timestamp 1640019720
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
<< locali >>
rect 59461 69615 59495 70193
rect 59553 70091 59587 70193
rect 88349 69955 88383 70125
rect 108313 69615 108347 69853
<<<<<<< HEAD
rect 204913 69683 204947 69921
rect 300869 69887 300903 70193
rect 209973 69071 210007 69717
rect 230489 69615 230523 69853
rect 301513 69343 301547 70193
rect 383853 69955 383887 70193
rect 388453 69683 388487 70261
rect 16865 3587 16899 3689
rect 43545 3315 43579 3689
rect 103805 3519 103839 4233
rect 103989 3451 104023 3961
rect 105645 3519 105679 3961
rect 399861 3961 400447 3995
rect 113833 3247 113867 3485
rect 116409 2907 116443 3417
=======
rect 204821 69683 204855 69921
rect 213469 69683 213503 69853
rect 296085 69819 296119 70261
rect 301513 69819 301547 70193
rect 214573 69275 214607 69649
rect 233801 69615 233835 69785
rect 301605 69343 301639 70193
rect 388545 69955 388579 70193
rect 388637 69343 388671 70193
rect 209973 69071 210007 69241
rect 16865 3587 16899 3689
rect 43545 3315 43579 3689
rect 106875 3485 107669 3519
rect 108313 3451 108347 3961
rect 399861 3961 400447 3995
rect 116409 2907 116443 3485
rect 116593 2975 116627 3417
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 160017 3383 160051 3689
rect 311357 3587 311391 3621
rect 311207 3553 311391 3587
rect 312587 3553 313289 3587
<<<<<<< HEAD
rect 316049 3451 316083 3689
rect 316141 3519 316175 3553
rect 316141 3485 316325 3519
rect 316049 3417 316233 3451
rect 337301 3315 337335 3825
rect 349445 3451 349479 3893
=======
rect 316141 3451 316175 3553
rect 337117 3043 337151 3757
rect 337301 3247 337335 3825
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 399861 3791 399895 3961
rect 400413 3927 400447 3961
rect 400321 3791 400355 3893
rect 400229 3519 400263 3757
<<<<<<< HEAD
rect 116593 2975 116627 3281
<< viali >>
rect 388453 70261 388487 70295
rect 59461 70193 59495 70227
rect 59553 70193 59587 70227
rect 300869 70193 300903 70227
rect 59553 70057 59587 70091
rect 88349 70125 88383 70159
rect 88349 69921 88383 69955
rect 204913 69921 204947 69955
rect 59461 69581 59495 69615
rect 108313 69853 108347 69887
rect 230489 69853 230523 69887
rect 300869 69853 300903 69887
rect 301513 70193 301547 70227
rect 204913 69649 204947 69683
rect 209973 69717 210007 69751
rect 108313 69581 108347 69615
rect 230489 69581 230523 69615
rect 383853 70193 383887 70227
rect 383853 69921 383887 69955
rect 388453 69649 388487 69683
rect 301513 69309 301547 69343
rect 209973 69037 210007 69071
rect 103805 4233 103839 4267
rect 16865 3689 16899 3723
rect 16865 3553 16899 3587
rect 43545 3689 43579 3723
rect 103805 3485 103839 3519
rect 103989 3961 104023 3995
rect 105645 3961 105679 3995
rect 349445 3893 349479 3927
rect 337301 3825 337335 3859
rect 160017 3689 160051 3723
rect 105645 3485 105679 3519
rect 113833 3485 113867 3519
rect 103989 3417 104023 3451
rect 43545 3281 43579 3315
rect 113833 3213 113867 3247
rect 116409 3417 116443 3451
rect 316049 3689 316083 3723
=======
rect 342269 2907 342303 3349
<< viali >>
rect 296085 70261 296119 70295
rect 59461 70193 59495 70227
rect 59553 70193 59587 70227
rect 59553 70057 59587 70091
rect 88349 70125 88383 70159
rect 88349 69921 88383 69955
rect 204821 69921 204855 69955
rect 59461 69581 59495 69615
rect 108313 69853 108347 69887
rect 204821 69649 204855 69683
rect 213469 69853 213503 69887
rect 233801 69785 233835 69819
rect 296085 69785 296119 69819
rect 301513 70193 301547 70227
rect 301513 69785 301547 69819
rect 301605 70193 301639 70227
rect 213469 69649 213503 69683
rect 214573 69649 214607 69683
rect 108313 69581 108347 69615
rect 233801 69581 233835 69615
rect 388545 70193 388579 70227
rect 388545 69921 388579 69955
rect 388637 70193 388671 70227
rect 301605 69309 301639 69343
rect 388637 69309 388671 69343
rect 209973 69241 210007 69275
rect 214573 69241 214607 69275
rect 209973 69037 210007 69071
rect 108313 3961 108347 3995
rect 16865 3689 16899 3723
rect 16865 3553 16899 3587
rect 43545 3689 43579 3723
rect 106841 3485 106875 3519
rect 107669 3485 107703 3519
rect 337301 3825 337335 3859
rect 337117 3757 337151 3791
rect 160017 3689 160051 3723
rect 108313 3417 108347 3451
rect 116409 3485 116443 3519
rect 43545 3281 43579 3315
rect 116593 3417 116627 3451
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 311357 3621 311391 3655
rect 311173 3553 311207 3587
rect 312553 3553 312587 3587
rect 313289 3553 313323 3587
rect 316141 3553 316175 3587
<<<<<<< HEAD
rect 316325 3485 316359 3519
rect 316233 3417 316267 3451
=======
rect 316141 3417 316175 3451
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 160017 3349 160051 3383
rect 400321 3893 400355 3927
rect 400413 3893 400447 3927
rect 399861 3757 399895 3791
rect 400229 3757 400263 3791
rect 400321 3757 400355 3791
rect 400229 3485 400263 3519
<<<<<<< HEAD
rect 349445 3417 349479 3451
rect 116593 3281 116627 3315
rect 337301 3281 337335 3315
rect 116593 2941 116627 2975
rect 116409 2873 116443 2907
=======
rect 337301 3213 337335 3247
rect 342269 3349 342303 3383
rect 337117 3009 337151 3043
rect 116593 2941 116627 2975
rect 116409 2873 116443 2907
rect 342269 2873 342303 2907
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
<< metal1 >>
rect 315942 700952 315948 701004
rect 316000 700992 316006 701004
rect 413646 700992 413652 701004
rect 316000 700964 413652 700992
rect 316000 700952 316006 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 325602 700884 325608 700936
rect 325660 700924 325666 700936
rect 429838 700924 429844 700936
rect 325660 700896 429844 700924
rect 325660 700884 325666 700896
rect 429838 700884 429844 700896
rect 429896 700884 429902 700936
rect 335262 700816 335268 700868
rect 335320 700856 335326 700868
rect 446122 700856 446128 700868
rect 335320 700828 446128 700856
rect 335320 700816 335326 700828
rect 446122 700816 446128 700828
rect 446180 700816 446186 700868
rect 346302 700748 346308 700800
rect 346360 700788 346366 700800
rect 462314 700788 462320 700800
rect 346360 700760 462320 700788
rect 346360 700748 346366 700760
rect 462314 700748 462320 700760
rect 462372 700748 462378 700800
rect 256602 700680 256608 700732
rect 256660 700720 256666 700732
rect 316310 700720 316316 700732
rect 256660 700692 316316 700720
rect 256660 700680 256666 700692
rect 316310 700680 316316 700692
rect 316368 700680 316374 700732
rect 355962 700680 355968 700732
rect 356020 700720 356026 700732
rect 478506 700720 478512 700732
rect 356020 700692 478512 700720
rect 356020 700680 356026 700692
rect 478506 700680 478512 700692
rect 478564 700680 478570 700732
rect 267550 700612 267556 700664
rect 267608 700652 267614 700664
rect 332502 700652 332508 700664
rect 267608 700624 332508 700652
rect 267608 700612 267614 700624
rect 332502 700612 332508 700624
rect 332560 700612 332566 700664
rect 365622 700612 365628 700664
rect 365680 700652 365686 700664
rect 494790 700652 494796 700664
rect 365680 700624 494796 700652
rect 365680 700612 365686 700624
rect 494790 700612 494796 700624
rect 494848 700612 494854 700664
rect 217962 700544 217968 700596
rect 218020 700584 218026 700596
rect 251450 700584 251456 700596
rect 218020 700556 251456 700584
rect 218020 700544 218026 700556
rect 251450 700544 251456 700556
rect 251508 700544 251514 700596
rect 277302 700544 277308 700596
rect 277360 700584 277366 700596
rect 348786 700584 348792 700596
rect 277360 700556 348792 700584
rect 277360 700544 277366 700556
rect 348786 700544 348792 700556
rect 348844 700544 348850 700596
rect 375282 700544 375288 700596
rect 375340 700584 375346 700596
rect 510982 700584 510988 700596
rect 375340 700556 510988 700584
rect 375340 700544 375346 700556
rect 510982 700544 510988 700556
rect 511040 700544 511046 700596
rect 227622 700476 227628 700528
rect 227680 700516 227686 700528
rect 267642 700516 267648 700528
rect 227680 700488 267648 700516
rect 227680 700476 227686 700488
rect 267642 700476 267648 700488
rect 267700 700476 267706 700528
rect 286962 700476 286968 700528
rect 287020 700516 287026 700528
rect 364978 700516 364984 700528
rect 287020 700488 364984 700516
rect 287020 700476 287026 700488
rect 364978 700476 364984 700488
rect 365036 700476 365042 700528
rect 384942 700476 384948 700528
rect 385000 700516 385006 700528
rect 527174 700516 527180 700528
rect 385000 700488 527180 700516
rect 385000 700476 385006 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 188982 700408 188988 700460
rect 189040 700448 189046 700460
rect 202782 700448 202788 700460
rect 189040 700420 202788 700448
rect 189040 700408 189046 700420
rect 202782 700408 202788 700420
rect 202840 700408 202846 700460
rect 237282 700408 237288 700460
rect 237340 700448 237346 700460
rect 283834 700448 283840 700460
rect 237340 700420 283840 700448
rect 237340 700408 237346 700420
rect 283834 700408 283840 700420
rect 283892 700408 283898 700460
rect 296622 700408 296628 700460
rect 296680 700448 296686 700460
rect 381170 700448 381176 700460
rect 296680 700420 381176 700448
rect 296680 700408 296686 700420
rect 381170 700408 381176 700420
rect 381228 700408 381234 700460
rect 394602 700408 394608 700460
rect 394660 700448 394666 700460
rect 543458 700448 543464 700460
rect 394660 700420 543464 700448
rect 394660 700408 394666 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 56778 700340 56784 700392
rect 56836 700380 56842 700392
rect 71038 700380 71044 700392
rect 56836 700352 71044 700380
rect 56836 700340 56842 700352
rect 71038 700340 71044 700352
rect 71096 700340 71102 700392
rect 177942 700340 177948 700392
rect 178000 700380 178006 700392
rect 186498 700380 186504 700392
rect 178000 700352 186504 700380
rect 178000 700340 178006 700352
rect 186498 700340 186504 700352
rect 186556 700340 186562 700392
rect 198642 700340 198648 700392
rect 198700 700380 198706 700392
rect 218974 700380 218980 700392
rect 198700 700352 218980 700380
rect 198700 700340 198706 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 220078 700340 220084 700392
rect 220136 700380 220142 700392
rect 235166 700380 235172 700392
rect 220136 700352 235172 700380
rect 220136 700340 220142 700352
rect 235166 700340 235172 700352
rect 235224 700340 235230 700392
rect 246942 700340 246948 700392
rect 247000 700380 247006 700392
rect 300118 700380 300124 700392
rect 247000 700352 300124 700380
rect 247000 700340 247006 700352
rect 300118 700340 300124 700352
rect 300176 700340 300182 700392
rect 306282 700340 306288 700392
rect 306340 700380 306346 700392
rect 397454 700380 397460 700392
rect 306340 700352 397460 700380
rect 306340 700340 306346 700352
rect 397454 700340 397460 700352
rect 397512 700340 397518 700392
rect 404262 700340 404268 700392
rect 404320 700380 404326 700392
rect 559650 700380 559656 700392
rect 404320 700352 559656 700380
rect 404320 700340 404326 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 62022 700272 62028 700324
rect 62080 700312 62086 700324
rect 575842 700312 575848 700324
rect 62080 700284 575848 700312
rect 62080 700272 62086 700284
rect 575842 700272 575848 700284
rect 575900 700272 575906 700324
rect 121638 700204 121644 700256
rect 121696 700244 121702 700256
rect 122742 700244 122748 700256
rect 121696 700216 122748 700244
rect 121696 700204 121702 700216
rect 122742 700204 122748 700216
rect 122800 700204 122806 700256
rect 154114 700068 154120 700120
rect 154172 700108 154178 700120
rect 155218 700108 155224 700120
rect 154172 700080 155224 700108
rect 154172 700068 154178 700080
rect 155218 700068 155224 700080
rect 155276 700068 155282 700120
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 169018 699660 169024 699712
rect 169076 699700 169082 699712
rect 170306 699700 170312 699712
rect 169076 699672 170312 699700
rect 169076 699660 169082 699672
rect 170306 699660 170312 699672
rect 170364 699660 170370 699712
rect 411898 696940 411904 696992
rect 411956 696980 411962 696992
rect 580166 696980 580172 696992
rect 411956 696952 580172 696980
rect 411956 696940 411962 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3142 683136 3148 683188
rect 3200 683176 3206 683188
rect 11698 683176 11704 683188
rect 3200 683148 11704 683176
rect 3200 683136 3206 683148
rect 11698 683136 11704 683148
rect 11756 683136 11762 683188
rect 406378 683136 406384 683188
rect 406436 683176 406442 683188
rect 580166 683176 580172 683188
rect 406436 683148 580172 683176
rect 406436 683136 406442 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 406470 670692 406476 670744
rect 406528 670732 406534 670744
rect 580166 670732 580172 670744
rect 406528 670704 580172 670732
rect 406528 670692 406534 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3142 656888 3148 656940
rect 3200 656928 3206 656940
rect 22738 656928 22744 656940
rect 3200 656900 22744 656928
rect 3200 656888 3206 656900
rect 22738 656888 22744 656900
rect 22796 656888 22802 656940
rect 410518 643084 410524 643136
rect 410576 643124 410582 643136
rect 580166 643124 580172 643136
rect 410576 643096 580172 643124
rect 410576 643084 410582 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3326 632068 3332 632120
rect 3384 632108 3390 632120
rect 14458 632108 14464 632120
rect 3384 632080 14464 632108
rect 3384 632068 3390 632080
rect 14458 632068 14464 632080
rect 14516 632068 14522 632120
rect 418798 630640 418804 630692
rect 418856 630680 418862 630692
rect 579982 630680 579988 630692
rect 418856 630652 579988 630680
rect 418856 630640 418862 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 2958 618264 2964 618316
rect 3016 618304 3022 618316
rect 35158 618304 35164 618316
rect 3016 618276 35164 618304
rect 3016 618264 3022 618276
rect 35158 618264 35164 618276
rect 35216 618264 35222 618316
rect 406562 616836 406568 616888
rect 406620 616876 406626 616888
rect 580166 616876 580172 616888
rect 406620 616848 580172 616876
rect 406620 616836 406626 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 25498 605860 25504 605872
rect 3384 605832 25504 605860
rect 3384 605820 3390 605832
rect 25498 605820 25504 605832
rect 25556 605820 25562 605872
rect 2774 592288 2780 592340
rect 2832 592328 2838 592340
rect 4798 592328 4804 592340
rect 2832 592300 4804 592328
rect 2832 592288 2838 592300
rect 4798 592288 4804 592300
rect 4856 592288 4862 592340
rect 406654 590656 406660 590708
rect 406712 590696 406718 590708
rect 579614 590696 579620 590708
rect 406712 590668 579620 590696
rect 406712 590656 406718 590668
rect 579614 590656 579620 590668
rect 579672 590656 579678 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 15838 579680 15844 579692
rect 3384 579652 15844 579680
rect 3384 579640 3390 579652
rect 15838 579640 15844 579652
rect 15896 579640 15902 579692
rect 406746 576852 406752 576904
rect 406804 576892 406810 576904
rect 579614 576892 579620 576904
rect 406804 576864 579620 576892
rect 406804 576852 406810 576864
rect 579614 576852 579620 576864
rect 579672 576852 579678 576904
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 36538 565876 36544 565888
rect 3108 565848 36544 565876
rect 3108 565836 3114 565848
rect 36538 565836 36544 565848
rect 36596 565836 36602 565888
rect 406838 563048 406844 563100
rect 406896 563088 406902 563100
rect 579890 563088 579896 563100
rect 406896 563060 579896 563088
rect 406896 563048 406902 563060
rect 579890 563048 579896 563060
rect 579948 563048 579954 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 29638 553432 29644 553444
rect 3384 553404 29644 553432
rect 3384 553392 3390 553404
rect 29638 553392 29644 553404
rect 29696 553392 29702 553444
rect 3326 539656 3332 539708
rect 3384 539696 3390 539708
rect 7558 539696 7564 539708
rect 3384 539668 7564 539696
rect 3384 539656 3390 539668
rect 7558 539656 7564 539668
rect 7616 539656 7622 539708
rect 407758 536800 407764 536852
rect 407816 536840 407822 536852
rect 580166 536840 580172 536852
rect 407816 536812 580172 536840
rect 407816 536800 407822 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3326 527144 3332 527196
rect 3384 527184 3390 527196
rect 17218 527184 17224 527196
rect 3384 527156 17224 527184
rect 3384 527144 3390 527156
rect 17218 527144 17224 527156
rect 17276 527144 17282 527196
rect 417418 524424 417424 524476
rect 417476 524464 417482 524476
rect 580166 524464 580172 524476
rect 417476 524436 580172 524464
rect 417476 524424 417482 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 32398 501004 32404 501016
rect 3292 500976 32404 501004
rect 3292 500964 3298 500976
rect 32398 500964 32404 500976
rect 32456 500964 32462 501016
rect 406930 484372 406936 484424
rect 406988 484412 406994 484424
rect 579614 484412 579620 484424
rect 406988 484384 579620 484412
rect 406988 484372 406994 484384
rect 579614 484372 579620 484384
rect 579672 484372 579678 484424
rect 2866 474716 2872 474768
rect 2924 474756 2930 474768
rect 18598 474756 18604 474768
rect 2924 474728 18604 474756
rect 2924 474716 2930 474728
rect 18598 474716 18604 474728
rect 18656 474716 18662 474768
rect 407022 470568 407028 470620
rect 407080 470608 407086 470620
rect 579982 470608 579988 470620
rect 407080 470580 579988 470608
rect 407080 470568 407086 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3050 462340 3056 462392
rect 3108 462380 3114 462392
rect 39298 462380 39304 462392
rect 3108 462352 39304 462380
rect 3108 462340 3114 462352
rect 39298 462340 39304 462352
rect 39356 462340 39362 462392
rect 2958 448536 2964 448588
rect 3016 448576 3022 448588
rect 33778 448576 33784 448588
rect 3016 448548 33784 448576
rect 3016 448536 3022 448548
rect 33778 448536 33784 448548
rect 33836 448536 33842 448588
rect 414658 430584 414664 430636
rect 414716 430624 414722 430636
rect 579982 430624 579988 430636
rect 414716 430596 579988 430624
rect 414716 430584 414722 430596
rect 579982 430584 579988 430596
rect 580040 430584 580046 430636
rect 2958 422288 2964 422340
rect 3016 422328 3022 422340
rect 21358 422328 21364 422340
rect 3016 422300 21364 422328
rect 3016 422288 3022 422300
rect 21358 422288 21364 422300
rect 21416 422288 21422 422340
rect 406286 418140 406292 418192
rect 406344 418180 406350 418192
rect 580166 418180 580172 418192
rect 406344 418152 580172 418180
rect 406344 418140 406350 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 406194 404336 406200 404388
rect 406252 404376 406258 404388
rect 580166 404376 580172 404388
rect 406252 404348 580172 404376
rect 406252 404336 406258 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 406102 378156 406108 378208
rect 406160 378196 406166 378208
rect 579798 378196 579804 378208
rect 406160 378168 579804 378196
rect 406160 378156 406166 378168
rect 579798 378156 579804 378168
rect 579856 378156 579862 378208
rect 60826 369792 60832 369844
rect 60884 369832 60890 369844
rect 62022 369832 62028 369844
rect 60884 369804 62028 369832
rect 60884 369792 60890 369804
rect 62022 369792 62028 369804
rect 62080 369792 62086 369844
rect 168098 369792 168104 369844
rect 168156 369832 168162 369844
rect 169018 369832 169024 369844
rect 168156 369804 169024 369832
rect 168156 369792 168162 369804
rect 169018 369792 169024 369804
rect 169076 369792 169082 369844
rect 217226 369792 217232 369844
rect 217284 369832 217290 369844
rect 217962 369832 217968 369844
rect 217284 369804 217968 369832
rect 217284 369792 217290 369804
rect 217962 369792 217968 369804
rect 218020 369792 218026 369844
rect 227070 369792 227076 369844
rect 227128 369832 227134 369844
rect 227622 369832 227628 369844
rect 227128 369804 227628 369832
rect 227128 369792 227134 369804
rect 227622 369792 227628 369804
rect 227680 369792 227686 369844
rect 286042 369792 286048 369844
rect 286100 369832 286106 369844
rect 286962 369832 286968 369844
rect 286100 369804 286968 369832
rect 286100 369792 286106 369804
rect 286962 369792 286968 369804
rect 287020 369792 287026 369844
rect 295886 369792 295892 369844
rect 295944 369832 295950 369844
rect 296622 369832 296628 369844
rect 295944 369804 296628 369832
rect 295944 369792 295950 369804
rect 296622 369792 296628 369804
rect 296680 369792 296686 369844
rect 305730 369792 305736 369844
rect 305788 369832 305794 369844
rect 306282 369832 306288 369844
rect 305788 369804 306288 369832
rect 305788 369792 305794 369804
rect 306282 369792 306288 369804
rect 306340 369792 306346 369844
rect 354858 369792 354864 369844
rect 354916 369832 354922 369844
rect 355962 369832 355968 369844
rect 354916 369804 355968 369832
rect 354916 369792 354922 369804
rect 355962 369792 355968 369804
rect 356020 369792 356026 369844
rect 364702 369792 364708 369844
rect 364760 369832 364766 369844
rect 365622 369832 365628 369844
rect 364760 369804 365628 369832
rect 364760 369792 364766 369804
rect 365622 369792 365628 369804
rect 365680 369792 365686 369844
rect 374546 369792 374552 369844
rect 374604 369832 374610 369844
rect 375282 369832 375288 369844
rect 374604 369804 375288 369832
rect 374604 369792 374610 369804
rect 375282 369792 375288 369804
rect 375340 369792 375346 369844
rect 384390 369792 384396 369844
rect 384448 369832 384454 369844
rect 384942 369832 384948 369844
rect 384448 369804 384948 369832
rect 384448 369792 384454 369804
rect 384942 369792 384948 369804
rect 385000 369792 385006 369844
rect 402974 369792 402980 369844
rect 403032 369832 403038 369844
rect 404262 369832 404268 369844
rect 403032 369804 404268 369832
rect 403032 369792 403038 369804
rect 404262 369792 404268 369804
rect 404320 369792 404326 369844
rect 197630 369656 197636 369708
rect 197688 369696 197694 369708
rect 198642 369696 198648 369708
rect 197688 369668 198648 369696
rect 197688 369656 197694 369668
rect 198642 369656 198648 369668
rect 198700 369656 198706 369708
rect 71038 369316 71044 369368
rect 71096 369356 71102 369368
rect 99282 369356 99288 369368
rect 71096 369328 99288 369356
rect 71096 369316 71102 369328
rect 99282 369316 99288 369328
rect 99340 369316 99346 369368
rect 41322 369248 41328 369300
rect 41380 369288 41386 369300
rect 89438 369288 89444 369300
rect 41380 369260 89444 369288
rect 41380 369248 41386 369260
rect 89438 369248 89444 369260
rect 89496 369248 89502 369300
rect 106182 369248 106188 369300
rect 106240 369288 106246 369300
rect 128814 369288 128820 369300
rect 106240 369260 128820 369288
rect 106240 369248 106246 369260
rect 128814 369248 128820 369260
rect 128872 369248 128878 369300
rect 24762 369180 24768 369232
rect 24820 369220 24826 369232
rect 79594 369220 79600 369232
rect 24820 369192 79600 369220
rect 24820 369180 24826 369192
rect 79594 369180 79600 369192
rect 79652 369180 79658 369232
rect 89622 369180 89628 369232
rect 89680 369220 89686 369232
rect 118970 369220 118976 369232
rect 89680 369192 118976 369220
rect 89680 369180 89686 369192
rect 118970 369180 118976 369192
rect 119028 369180 119034 369232
rect 137922 369180 137928 369232
rect 137980 369220 137986 369232
rect 148410 369220 148416 369232
rect 137980 369192 148416 369220
rect 137980 369180 137986 369192
rect 148410 369180 148416 369192
rect 148468 369180 148474 369232
rect 155218 369180 155224 369232
rect 155276 369220 155282 369232
rect 158254 369220 158260 369232
rect 155276 369192 158260 369220
rect 155276 369180 155282 369192
rect 158254 369180 158260 369192
rect 158312 369180 158318 369232
rect 8202 369112 8208 369164
rect 8260 369152 8266 369164
rect 69750 369152 69756 369164
rect 8260 369124 69756 369152
rect 8260 369112 8266 369124
rect 69750 369112 69756 369124
rect 69808 369112 69814 369164
rect 73062 369112 73068 369164
rect 73120 369152 73126 369164
rect 109126 369152 109132 369164
rect 73120 369124 109132 369152
rect 73120 369112 73126 369124
rect 109126 369112 109132 369124
rect 109184 369112 109190 369164
rect 122742 369112 122748 369164
rect 122800 369152 122806 369164
rect 138566 369152 138572 369164
rect 122800 369124 138572 369152
rect 122800 369112 122806 369124
rect 138566 369112 138572 369124
rect 138624 369112 138630 369164
rect 187786 369112 187792 369164
rect 187844 369152 187850 369164
rect 188982 369152 188988 369164
rect 187844 369124 188988 369152
rect 187844 369112 187850 369124
rect 188982 369112 188988 369124
rect 189040 369112 189046 369164
rect 207474 369112 207480 369164
rect 207532 369152 207538 369164
rect 220078 369152 220084 369164
rect 207532 369124 220084 369152
rect 207532 369112 207538 369124
rect 220078 369112 220084 369124
rect 220136 369112 220142 369164
rect 345106 369112 345112 369164
rect 345164 369152 345170 369164
rect 346302 369152 346308 369164
rect 345164 369124 346308 369152
rect 345164 369112 345170 369124
rect 346302 369112 346308 369124
rect 346360 369112 346366 369164
rect 266446 369044 266452 369096
rect 266504 369084 266510 369096
rect 267642 369084 267648 369096
rect 266504 369056 267648 369084
rect 266504 369044 266510 369056
rect 267642 369044 267648 369056
rect 267700 369044 267706 369096
rect 276290 368976 276296 369028
rect 276348 369016 276354 369028
rect 277302 369016 277308 369028
rect 276348 368988 277308 369016
rect 276348 368976 276354 368988
rect 277302 368976 277308 368988
rect 277360 368976 277366 369028
rect 3418 365644 3424 365696
rect 3476 365684 3482 365696
rect 57422 365684 57428 365696
rect 3476 365656 57428 365684
rect 3476 365644 3482 365656
rect 57422 365644 57428 365656
rect 57480 365644 57486 365696
rect 406010 364964 406016 365016
rect 406068 365004 406074 365016
rect 411898 365004 411904 365016
rect 406068 364976 411904 365004
rect 406068 364964 406074 364976
rect 411898 364964 411904 364976
rect 411956 364964 411962 365016
rect 411990 364352 411996 364404
rect 412048 364392 412054 364404
rect 580166 364392 580172 364404
rect 412048 364364 580172 364392
rect 412048 364352 412054 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 11698 361496 11704 361548
rect 11756 361536 11762 361548
rect 57146 361536 57152 361548
rect 11756 361508 57152 361536
rect 11756 361496 11762 361508
rect 57146 361496 57152 361508
rect 57204 361496 57210 361548
rect 3510 355988 3516 356040
rect 3568 356028 3574 356040
rect 57238 356028 57244 356040
rect 3568 356000 57244 356028
rect 3568 355988 3574 356000
rect 57238 355988 57244 356000
rect 57296 355988 57302 356040
rect 406378 351908 406384 351960
rect 406436 351948 406442 351960
rect 580166 351948 580172 351960
rect 406436 351920 580172 351948
rect 406436 351908 406442 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 22738 350480 22744 350532
rect 22796 350520 22802 350532
rect 57606 350520 57612 350532
rect 22796 350492 57612 350520
rect 22796 350480 22802 350492
rect 57606 350480 57612 350492
rect 57664 350480 57670 350532
rect 406470 349052 406476 349104
rect 406528 349092 406534 349104
rect 580074 349092 580080 349104
rect 406528 349064 580080 349092
rect 406528 349052 406534 349064
rect 580074 349052 580080 349064
rect 580132 349052 580138 349104
rect 3602 344972 3608 345024
rect 3660 345012 3666 345024
rect 57606 345012 57612 345024
rect 3660 344984 57612 345012
rect 3660 344972 3666 344984
rect 57606 344972 57612 344984
rect 57664 344972 57670 345024
rect 406470 343340 406476 343392
rect 406528 343380 406534 343392
rect 410518 343380 410524 343392
rect 406528 343352 410524 343380
rect 406528 343340 406534 343352
rect 410518 343340 410524 343352
rect 410576 343340 410582 343392
rect 14458 339396 14464 339448
rect 14516 339436 14522 339448
rect 57606 339436 57612 339448
rect 14516 339408 57612 339436
rect 14516 339396 14522 339408
rect 57606 339396 57612 339408
rect 57664 339396 57670 339448
rect 406470 338036 406476 338088
rect 406528 338076 406534 338088
rect 418798 338076 418804 338088
rect 406528 338048 418804 338076
rect 406528 338036 406534 338048
rect 418798 338036 418804 338048
rect 418856 338036 418862 338088
rect 35158 333888 35164 333940
rect 35216 333928 35222 333940
rect 57606 333928 57612 333940
rect 35216 333900 57612 333928
rect 35216 333888 35222 333900
rect 57606 333888 57612 333900
rect 57664 333888 57670 333940
rect 25498 328380 25504 328432
rect 25556 328420 25562 328432
rect 57330 328420 57336 328432
rect 25556 328392 57336 328420
rect 25556 328380 25562 328392
rect 57330 328380 57336 328392
rect 57388 328380 57394 328432
rect 406562 327020 406568 327072
rect 406620 327060 406626 327072
rect 580350 327060 580356 327072
rect 406620 327032 580356 327060
rect 406620 327020 406626 327032
rect 580350 327020 580356 327032
rect 580408 327020 580414 327072
rect 406470 324300 406476 324352
rect 406528 324340 406534 324352
rect 580166 324340 580172 324352
rect 406528 324312 580172 324340
rect 406528 324300 406534 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 4798 322872 4804 322924
rect 4856 322912 4862 322924
rect 57330 322912 57336 322924
rect 4856 322884 57336 322912
rect 4856 322872 4862 322884
rect 57330 322872 57336 322884
rect 57388 322872 57394 322924
rect 15838 317364 15844 317416
rect 15896 317404 15902 317416
rect 57606 317404 57612 317416
rect 15896 317376 57612 317404
rect 15896 317364 15902 317376
rect 57606 317364 57612 317376
rect 57664 317364 57670 317416
rect 406562 311856 406568 311908
rect 406620 311896 406626 311908
rect 580166 311896 580172 311908
rect 406620 311868 580172 311896
rect 406620 311856 406626 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 36538 310428 36544 310480
rect 36596 310468 36602 310480
rect 57606 310468 57612 310480
rect 36596 310440 57612 310468
rect 36596 310428 36602 310440
rect 57606 310428 57612 310440
rect 57664 310428 57670 310480
rect 29638 304920 29644 304972
rect 29696 304960 29702 304972
rect 57422 304960 57428 304972
rect 29696 304932 57428 304960
rect 29696 304920 29702 304932
rect 57422 304920 57428 304932
rect 57480 304920 57486 304972
rect 406838 304920 406844 304972
rect 406896 304960 406902 304972
rect 580442 304960 580448 304972
rect 406896 304932 580448 304960
rect 406896 304920 406902 304932
rect 580442 304920 580448 304932
rect 580500 304920 580506 304972
rect 7558 299412 7564 299464
rect 7616 299452 7622 299464
rect 57606 299452 57612 299464
rect 7616 299424 57612 299452
rect 7616 299412 7622 299424
rect 57606 299412 57612 299424
rect 57664 299412 57670 299464
rect 405826 299276 405832 299328
rect 405884 299316 405890 299328
rect 407758 299316 407764 299328
rect 405884 299288 407764 299316
rect 405884 299276 405890 299288
rect 407758 299276 407764 299288
rect 407816 299276 407822 299328
rect 406654 298120 406660 298172
rect 406712 298160 406718 298172
rect 580166 298160 580172 298172
rect 406712 298132 580172 298160
rect 406712 298120 406718 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 17218 293904 17224 293956
rect 17276 293944 17282 293956
rect 57606 293944 57612 293956
rect 17276 293916 57612 293944
rect 17276 293904 17282 293916
rect 57606 293904 57612 293916
rect 57664 293904 57670 293956
rect 406838 292476 406844 292528
rect 406896 292516 406902 292528
rect 417418 292516 417424 292528
rect 406896 292488 417424 292516
rect 406896 292476 406902 292488
rect 417418 292476 417424 292488
rect 417476 292476 417482 292528
rect 3694 288328 3700 288380
rect 3752 288368 3758 288380
rect 57606 288368 57612 288380
rect 3752 288340 57612 288368
rect 3752 288328 3758 288340
rect 57606 288328 57612 288340
rect 57664 288328 57670 288380
rect 406838 286968 406844 287020
rect 406896 287008 406902 287020
rect 580534 287008 580540 287020
rect 406896 286980 580540 287008
rect 406896 286968 406902 286980
rect 580534 286968 580540 286980
rect 580592 286968 580598 287020
rect 32398 282820 32404 282872
rect 32456 282860 32462 282872
rect 57606 282860 57612 282872
rect 32456 282832 57612 282860
rect 32456 282820 32462 282832
rect 57606 282820 57612 282832
rect 57664 282820 57670 282872
rect 406838 281460 406844 281512
rect 406896 281500 406902 281512
rect 580626 281500 580632 281512
rect 406896 281472 580632 281500
rect 406896 281460 406902 281472
rect 580626 281460 580632 281472
rect 580684 281460 580690 281512
rect 3786 277312 3792 277364
rect 3844 277352 3850 277364
rect 57606 277352 57612 277364
rect 3844 277324 57612 277352
rect 3844 277312 3850 277324
rect 57606 277312 57612 277324
rect 57664 277312 57670 277364
rect 406746 271872 406752 271924
rect 406804 271912 406810 271924
rect 580166 271912 580172 271924
rect 406804 271884 580172 271912
rect 406804 271872 406810 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 18598 271804 18604 271856
rect 18656 271844 18662 271856
rect 57514 271844 57520 271856
rect 18656 271816 57520 271844
rect 18656 271804 18662 271816
rect 57514 271804 57520 271816
rect 57572 271804 57578 271856
rect 39298 266296 39304 266348
rect 39356 266336 39362 266348
rect 57330 266336 57336 266348
rect 39356 266308 57336 266336
rect 39356 266296 39362 266308
rect 57330 266296 57336 266308
rect 57388 266296 57394 266348
rect 407022 264868 407028 264920
rect 407080 264908 407086 264920
rect 580718 264908 580724 264920
rect 407080 264880 580724 264908
rect 407080 264868 407086 264880
rect 580718 264868 580724 264880
rect 580776 264868 580782 264920
rect 33778 260788 33784 260840
rect 33836 260828 33842 260840
rect 57422 260828 57428 260840
rect 33836 260800 57428 260828
rect 33836 260788 33842 260800
rect 57422 260788 57428 260800
rect 57480 260788 57486 260840
rect 406930 259360 406936 259412
rect 406988 259400 406994 259412
rect 580810 259400 580816 259412
rect 406988 259372 580816 259400
rect 406988 259360 406994 259372
rect 580810 259360 580816 259372
rect 580868 259360 580874 259412
rect 406838 258068 406844 258120
rect 406896 258108 406902 258120
rect 580166 258108 580172 258120
rect 406896 258080 580172 258108
rect 406896 258068 406902 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 3878 255212 3884 255264
rect 3936 255252 3942 255264
rect 57606 255252 57612 255264
rect 3936 255224 57612 255252
rect 3936 255212 3942 255224
rect 57606 255212 57612 255224
rect 57664 255212 57670 255264
rect 407022 252832 407028 252884
rect 407080 252872 407086 252884
rect 414658 252872 414664 252884
rect 407080 252844 414664 252872
rect 407080 252832 407086 252844
rect 414658 252832 414664 252844
rect 414716 252832 414722 252884
rect 21358 249704 21364 249756
rect 21416 249744 21422 249756
rect 57238 249744 57244 249756
rect 21416 249716 57244 249744
rect 21416 249704 21422 249716
rect 57238 249704 57244 249716
rect 57296 249704 57302 249756
rect 406930 244264 406936 244316
rect 406988 244304 406994 244316
rect 580166 244304 580172 244316
rect 406988 244276 580172 244304
rect 406988 244264 406994 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 3970 244196 3976 244248
rect 4028 244236 4034 244248
rect 57422 244236 57428 244248
rect 4028 244208 57428 244236
rect 4028 244196 4034 244208
rect 57422 244196 57428 244208
rect 57480 244196 57486 244248
rect 4062 238688 4068 238740
rect 4120 238728 4126 238740
rect 57606 238728 57612 238740
rect 4120 238700 57612 238728
rect 4120 238688 4126 238700
rect 57606 238688 57612 238700
rect 57664 238688 57670 238740
rect 407022 235900 407028 235952
rect 407080 235940 407086 235952
rect 580902 235940 580908 235952
rect 407080 235912 580908 235940
rect 407080 235900 407086 235912
rect 580902 235900 580908 235912
rect 580960 235900 580966 235952
rect 3326 233180 3332 233232
rect 3384 233220 3390 233232
rect 57606 233220 57612 233232
rect 3384 233192 57612 233220
rect 3384 233180 3390 233192
rect 57606 233180 57612 233192
rect 57664 233180 57670 233232
rect 407022 231820 407028 231872
rect 407080 231860 407086 231872
rect 579614 231860 579620 231872
rect 407080 231832 579620 231860
rect 407080 231820 407086 231832
rect 579614 231820 579620 231832
rect 579672 231820 579678 231872
rect 3234 227672 3240 227724
rect 3292 227712 3298 227724
rect 57606 227712 57612 227724
rect 3292 227684 57612 227712
rect 3292 227672 3298 227684
rect 57606 227672 57612 227684
rect 57664 227672 57670 227724
rect 406286 224612 406292 224664
rect 406344 224652 406350 224664
rect 411990 224652 411996 224664
rect 406344 224624 411996 224652
rect 406344 224612 406350 224624
rect 411990 224612 411996 224624
rect 412048 224612 412054 224664
rect 3418 222096 3424 222148
rect 3476 222136 3482 222148
rect 57606 222136 57612 222148
rect 3476 222108 57612 222136
rect 3476 222096 3482 222108
rect 57606 222096 57612 222108
rect 57664 222096 57670 222148
rect 406286 218016 406292 218068
rect 406344 218056 406350 218068
rect 580166 218056 580172 218068
rect 406344 218028 580172 218056
rect 406344 218016 406350 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 3510 216588 3516 216640
rect 3568 216628 3574 216640
rect 57054 216628 57060 216640
rect 3568 216600 57060 216628
rect 3568 216588 3574 216600
rect 57054 216588 57060 216600
rect 57112 216588 57118 216640
rect 406378 213868 406384 213920
rect 406436 213908 406442 213920
rect 580258 213908 580264 213920
rect 406436 213880 580264 213908
rect 406436 213868 406442 213880
rect 580258 213868 580264 213880
rect 580316 213868 580322 213920
rect 3602 211080 3608 211132
rect 3660 211120 3666 211132
rect 56778 211120 56784 211132
rect 3660 211092 56784 211120
rect 3660 211080 3666 211092
rect 56778 211080 56784 211092
rect 56836 211080 56842 211132
rect 406378 205640 406384 205692
rect 406436 205680 406442 205692
rect 580166 205680 580172 205692
rect 406436 205652 580172 205680
rect 406436 205640 406442 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 3142 205572 3148 205624
rect 3200 205612 3206 205624
rect 57606 205612 57612 205624
rect 3200 205584 57612 205612
rect 3200 205572 3206 205584
rect 57606 205572 57612 205584
rect 57664 205572 57670 205624
rect 3050 200064 3056 200116
rect 3108 200104 3114 200116
rect 57606 200104 57612 200116
rect 3108 200076 57612 200104
rect 3108 200064 3114 200076
rect 57606 200064 57612 200076
rect 57664 200064 57670 200116
rect 2958 194488 2964 194540
rect 3016 194528 3022 194540
rect 57606 194528 57612 194540
rect 3016 194500 57612 194528
rect 3016 194488 3022 194500
rect 57606 194488 57612 194500
rect 57664 194488 57670 194540
rect 406470 191836 406476 191888
rect 406528 191876 406534 191888
rect 580166 191876 580172 191888
rect 406528 191848 580172 191876
rect 406528 191836 406534 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 406746 191768 406752 191820
rect 406804 191808 406810 191820
rect 580350 191808 580356 191820
rect 406804 191780 580356 191808
rect 406804 191768 406810 191780
rect 580350 191768 580356 191780
rect 580408 191768 580414 191820
rect 3694 188980 3700 189032
rect 3752 189020 3758 189032
rect 57606 189020 57612 189032
rect 3752 188992 57612 189020
rect 3752 188980 3758 188992
rect 57606 188980 57612 188992
rect 57664 188980 57670 189032
rect 3786 183472 3792 183524
rect 3844 183512 3850 183524
rect 57606 183512 57612 183524
rect 3844 183484 57612 183512
rect 3844 183472 3850 183484
rect 57606 183472 57612 183484
rect 57664 183472 57670 183524
rect 406562 178032 406568 178084
rect 406620 178072 406626 178084
rect 580166 178072 580172 178084
rect 406620 178044 580172 178072
rect 406620 178032 406626 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 2866 177964 2872 178016
rect 2924 178004 2930 178016
rect 56686 178004 56692 178016
rect 2924 177976 56692 178004
rect 2924 177964 2930 177976
rect 56686 177964 56692 177976
rect 56744 177964 56750 178016
rect 3878 172456 3884 172508
rect 3936 172496 3942 172508
rect 57606 172496 57612 172508
rect 3936 172468 57612 172496
rect 3936 172456 3942 172468
rect 57606 172456 57612 172468
rect 57664 172456 57670 172508
rect 3970 166948 3976 167000
rect 4028 166988 4034 167000
rect 57606 166988 57612 167000
rect 4028 166960 57612 166988
rect 4028 166948 4034 166960
rect 57606 166948 57612 166960
rect 57664 166948 57670 167000
rect 406654 165588 406660 165640
rect 406712 165628 406718 165640
rect 580166 165628 580172 165640
rect 406712 165600 580172 165628
rect 406712 165588 406718 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 3418 161372 3424 161424
rect 3476 161412 3482 161424
rect 57606 161412 57612 161424
rect 3476 161384 57612 161412
rect 3476 161372 3482 161384
rect 57606 161372 57612 161384
rect 57664 161372 57670 161424
rect 3510 155864 3516 155916
rect 3568 155904 3574 155916
rect 57606 155904 57612 155916
rect 3568 155876 57612 155904
rect 3568 155864 3574 155876
rect 57606 155864 57612 155876
rect 57664 155864 57670 155916
rect 406378 151784 406384 151836
rect 406436 151824 406442 151836
rect 579982 151824 579988 151836
rect 406436 151796 579988 151824
rect 406436 151784 406442 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 3602 150356 3608 150408
rect 3660 150396 3666 150408
rect 56870 150396 56876 150408
rect 3660 150368 56876 150396
rect 3660 150356 3666 150368
rect 56870 150356 56876 150368
rect 56928 150356 56934 150408
rect 3694 144848 3700 144900
rect 3752 144888 3758 144900
rect 57514 144888 57520 144900
rect 3752 144860 57520 144888
rect 3752 144848 3758 144860
rect 57514 144848 57520 144860
rect 57572 144848 57578 144900
rect 3786 139340 3792 139392
rect 3844 139380 3850 139392
rect 57514 139380 57520 139392
rect 3844 139352 57520 139380
rect 3844 139340 3850 139352
rect 57514 139340 57520 139352
rect 57572 139340 57578 139392
rect 406470 137980 406476 138032
rect 406528 138020 406534 138032
rect 580166 138020 580172 138032
rect 406528 137992 580172 138020
rect 406528 137980 406534 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 3418 133832 3424 133884
rect 3476 133872 3482 133884
rect 57514 133872 57520 133884
rect 3476 133844 57520 133872
rect 3476 133832 3482 133844
rect 57514 133832 57520 133844
rect 57572 133832 57578 133884
rect 3510 128256 3516 128308
rect 3568 128296 3574 128308
rect 56962 128296 56968 128308
rect 3568 128268 56968 128296
rect 3568 128256 3574 128268
rect 56962 128256 56968 128268
rect 57020 128256 57026 128308
rect 407022 125604 407028 125656
rect 407080 125644 407086 125656
rect 580166 125644 580172 125656
rect 407080 125616 580172 125644
rect 407080 125604 407086 125616
rect 580166 125604 580172 125616
rect 580224 125604 580230 125656
rect 3602 122748 3608 122800
rect 3660 122788 3666 122800
rect 57054 122788 57060 122800
rect 3660 122760 57060 122788
rect 3660 122748 3666 122760
rect 57054 122748 57060 122760
rect 57112 122748 57118 122800
rect 3418 115948 3424 116000
rect 3476 115988 3482 116000
rect 57606 115988 57612 116000
rect 3476 115960 57612 115988
rect 3476 115948 3482 115960
rect 57606 115948 57612 115960
rect 57664 115948 57670 116000
rect 406378 113092 406384 113144
rect 406436 113132 406442 113144
rect 579798 113132 579804 113144
rect 406436 113104 579804 113132
rect 406436 113092 406442 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3510 110440 3516 110492
rect 3568 110480 3574 110492
rect 57606 110480 57612 110492
rect 3568 110452 57612 110480
rect 3568 110440 3574 110452
rect 57606 110440 57612 110452
rect 57664 110440 57670 110492
rect 3418 104864 3424 104916
rect 3476 104904 3482 104916
rect 57422 104904 57428 104916
rect 3476 104876 57428 104904
rect 3476 104864 3482 104876
rect 57422 104864 57428 104876
rect 57480 104864 57486 104916
rect 406470 100648 406476 100700
rect 406528 100688 406534 100700
rect 580166 100688 580172 100700
rect 406528 100660 580172 100688
rect 406528 100648 406534 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3878 99356 3884 99408
rect 3936 99396 3942 99408
rect 57422 99396 57428 99408
rect 3936 99368 57428 99396
rect 3936 99356 3942 99368
rect 57422 99356 57428 99368
rect 57480 99356 57486 99408
rect 3786 93848 3792 93900
rect 3844 93888 3850 93900
rect 57606 93888 57612 93900
rect 3844 93860 57612 93888
rect 3844 93848 3850 93860
rect 57606 93848 57612 93860
rect 57664 93848 57670 93900
rect 3694 88340 3700 88392
rect 3752 88380 3758 88392
rect 57514 88380 57520 88392
rect 3752 88352 57520 88380
rect 3752 88340 3758 88352
rect 57514 88340 57520 88352
rect 57572 88340 57578 88392
rect 406378 86912 406384 86964
rect 406436 86952 406442 86964
rect 580166 86952 580172 86964
rect 406436 86924 580172 86952
rect 406436 86912 406442 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3602 82832 3608 82884
rect 3660 82872 3666 82884
rect 57422 82872 57428 82884
rect 3660 82844 57428 82872
rect 3660 82832 3666 82844
rect 57422 82832 57428 82844
rect 57480 82832 57486 82884
rect 3510 77256 3516 77308
rect 3568 77296 3574 77308
rect 57514 77296 57520 77308
rect 3568 77268 57520 77296
rect 3568 77256 3574 77268
rect 57514 77256 57520 77268
rect 57572 77256 57578 77308
rect 406838 73108 406844 73160
rect 406896 73148 406902 73160
rect 580166 73148 580172 73160
rect 406896 73120 580172 73148
rect 406896 73108 406902 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3418 71748 3424 71800
rect 3476 71788 3482 71800
rect 57422 71788 57428 71800
rect 3476 71760 57428 71788
rect 3476 71748 3482 71760
rect 57422 71748 57428 71760
rect 57480 71748 57486 71800
rect 60826 71748 60832 71800
rect 60884 71788 60890 71800
rect 62061 71788 62067 71800
rect 60884 71760 62067 71788
rect 60884 71748 60890 71760
rect 62061 71748 62067 71760
rect 62119 71748 62125 71800
rect 97994 71748 98000 71800
rect 98052 71788 98058 71800
rect 99045 71788 99051 71800
rect 98052 71760 99051 71788
rect 98052 71748 98058 71760
rect 99045 71748 99051 71760
rect 99103 71748 99109 71800
rect 100754 71748 100760 71800
rect 100812 71788 100818 71800
rect 101836 71788 101842 71800
rect 100812 71760 101842 71788
rect 100812 71748 100818 71760
rect 101836 71748 101842 71760
rect 101894 71748 101900 71800
rect 109126 71748 109132 71800
rect 109184 71788 109190 71800
rect 110210 71788 110216 71800
rect 109184 71760 110216 71788
rect 109184 71748 109190 71760
rect 110210 71748 110216 71760
rect 110268 71748 110274 71800
rect 114554 71748 114560 71800
rect 114612 71788 114618 71800
rect 115792 71788 115798 71800
rect 114612 71760 115798 71788
rect 114612 71748 114618 71760
rect 115792 71748 115798 71760
rect 115850 71748 115856 71800
rect 116026 71748 116032 71800
rect 116084 71788 116090 71800
rect 117188 71788 117194 71800
rect 116084 71760 117194 71788
rect 116084 71748 116090 71760
rect 117188 71748 117194 71760
rect 117246 71748 117252 71800
rect 117314 71748 117320 71800
rect 117372 71788 117378 71800
rect 118583 71788 118589 71800
rect 117372 71760 118589 71788
rect 117372 71748 117378 71760
rect 118583 71748 118589 71760
rect 118641 71748 118647 71800
rect 118786 71748 118792 71800
rect 118844 71788 118850 71800
rect 119979 71788 119985 71800
rect 118844 71760 119985 71788
rect 118844 71748 118850 71760
rect 119979 71748 119985 71760
rect 120037 71748 120043 71800
rect 120166 71748 120172 71800
rect 120224 71788 120230 71800
rect 121374 71788 121380 71800
rect 120224 71760 121380 71788
rect 120224 71748 120230 71760
rect 121374 71748 121380 71760
rect 121432 71748 121438 71800
rect 230474 71748 230480 71800
rect 230532 71788 230538 71800
rect 231627 71788 231633 71800
rect 230532 71760 231633 71788
rect 230532 71748 230538 71760
rect 231627 71748 231633 71760
rect 231685 71748 231691 71800
rect 234706 71748 234712 71800
rect 234764 71788 234770 71800
rect 235814 71788 235820 71800
rect 234764 71760 235820 71788
rect 234764 71748 234770 71760
rect 235814 71748 235820 71760
rect 235872 71748 235878 71800
rect 236086 71748 236092 71800
rect 236144 71788 236150 71800
rect 237209 71788 237215 71800
rect 236144 71760 237215 71788
rect 236144 71748 236150 71760
rect 237209 71748 237215 71760
rect 237267 71748 237273 71800
rect 237374 71748 237380 71800
rect 237432 71788 237438 71800
rect 238605 71788 238611 71800
rect 237432 71760 238611 71788
rect 237432 71748 237438 71760
rect 238605 71748 238611 71760
rect 238663 71748 238669 71800
rect 240134 71748 240140 71800
rect 240192 71788 240198 71800
rect 241396 71788 241402 71800
rect 240192 71760 241402 71788
rect 240192 71748 240198 71760
rect 241396 71748 241402 71760
rect 241454 71748 241460 71800
rect 321554 71748 321560 71800
rect 321612 71788 321618 71800
rect 322341 71788 322347 71800
rect 321612 71760 322347 71788
rect 321612 71748 321618 71760
rect 322341 71748 322347 71760
rect 322399 71748 322405 71800
rect 324314 71748 324320 71800
rect 324372 71788 324378 71800
rect 325132 71788 325138 71800
rect 324372 71760 325138 71788
rect 324372 71748 324378 71760
rect 325132 71748 325138 71760
rect 325190 71748 325196 71800
rect 327074 71748 327080 71800
rect 327132 71788 327138 71800
rect 327923 71788 327929 71800
rect 327132 71760 327929 71788
rect 327132 71748 327138 71760
rect 327923 71748 327929 71760
rect 327981 71748 327987 71800
rect 328454 71748 328460 71800
rect 328512 71788 328518 71800
rect 329319 71788 329325 71800
rect 328512 71760 329325 71788
rect 328512 71748 328518 71760
rect 329319 71748 329325 71760
rect 329377 71748 329383 71800
rect 329834 71748 329840 71800
rect 329892 71788 329898 71800
rect 330714 71788 330720 71800
rect 329892 71760 330720 71788
rect 329892 71748 329898 71760
rect 330714 71748 330720 71760
rect 330772 71748 330778 71800
rect 331214 71748 331220 71800
rect 331272 71788 331278 71800
rect 332110 71788 332116 71800
rect 331272 71760 332116 71788
rect 331272 71748 331278 71760
rect 332110 71748 332116 71760
rect 332168 71748 332174 71800
rect 333974 71748 333980 71800
rect 334032 71788 334038 71800
rect 334901 71788 334907 71800
rect 334032 71760 334907 71788
rect 334032 71748 334038 71760
rect 334901 71748 334907 71760
rect 334959 71748 334965 71800
rect 335446 71748 335452 71800
rect 335504 71788 335510 71800
rect 336297 71788 336303 71800
rect 335504 71760 336303 71788
rect 335504 71748 335510 71760
rect 336297 71748 336303 71760
rect 336355 71748 336361 71800
rect 338114 71748 338120 71800
rect 338172 71788 338178 71800
rect 339088 71788 339094 71800
rect 338172 71760 339094 71788
rect 338172 71748 338178 71760
rect 339088 71748 339094 71760
rect 339146 71748 339152 71800
rect 340966 71748 340972 71800
rect 341024 71788 341030 71800
rect 341879 71788 341885 71800
rect 341024 71760 341885 71788
rect 341024 71748 341030 71760
rect 341879 71748 341885 71760
rect 341937 71748 341943 71800
rect 349246 71748 349252 71800
rect 349304 71788 349310 71800
rect 350253 71788 350259 71800
rect 349304 71760 350259 71788
rect 349304 71748 349310 71760
rect 350253 71748 350259 71760
rect 350311 71748 350317 71800
rect 53098 70320 53104 70372
rect 53156 70360 53162 70372
rect 64138 70360 64144 70372
rect 53156 70332 64144 70360
rect 53156 70320 53162 70332
rect 64138 70320 64144 70332
rect 64196 70320 64202 70372
rect 148962 70320 148968 70372
rect 149020 70360 149026 70372
rect 227438 70360 227444 70372
rect 149020 70332 227444 70360
rect 149020 70320 149026 70332
rect 227438 70320 227444 70332
rect 227496 70320 227502 70372
rect 265802 70320 265808 70372
rect 265860 70360 265866 70372
<<<<<<< HEAD
rect 295978 70360 295984 70372
rect 265860 70332 295984 70360
rect 265860 70320 265866 70332
rect 295978 70320 295984 70332
rect 296036 70320 296042 70372
=======
rect 295886 70360 295892 70372
rect 265860 70332 295892 70360
rect 265860 70320 265866 70332
rect 295886 70320 295892 70332
rect 295944 70320 295950 70372
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 299382 70320 299388 70372
rect 299440 70360 299446 70372
rect 346026 70360 346032 70372
rect 299440 70332 346032 70360
rect 299440 70320 299446 70332
rect 346026 70320 346032 70332
rect 346084 70320 346090 70372
<<<<<<< HEAD
rect 375374 70320 375380 70372
rect 375432 70360 375438 70372
rect 447134 70360 447140 70372
rect 375432 70332 447140 70360
rect 375432 70320 375438 70332
rect 447134 70320 447140 70332
rect 447192 70320 447198 70372
=======
rect 373994 70320 374000 70372
rect 374052 70360 374058 70372
rect 440234 70360 440240 70372
rect 374052 70332 440240 70360
rect 374052 70320 374058 70332
rect 440234 70320 440240 70332
rect 440292 70320 440298 70372
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 41322 70252 41328 70304
rect 41380 70292 41386 70304
rect 67634 70292 67640 70304
rect 41380 70264 67640 70292
rect 41380 70252 41386 70264
rect 67634 70252 67640 70264
rect 67692 70252 67698 70304
rect 121362 70252 121368 70304
rect 121420 70292 121426 70304
rect 128354 70292 128360 70304
rect 121420 70264 128360 70292
rect 121420 70252 121426 70264
rect 128354 70252 128360 70264
rect 128412 70252 128418 70304
rect 141970 70252 141976 70304
rect 142028 70292 142034 70304
rect 226058 70292 226064 70304
rect 142028 70264 226064 70292
rect 142028 70252 142034 70264
rect 226058 70252 226064 70264
rect 226116 70252 226122 70304
<<<<<<< HEAD
rect 287698 70252 287704 70304
rect 287756 70292 287762 70304
rect 325786 70292 325792 70304
rect 287756 70264 325792 70292
rect 287756 70252 287762 70264
=======
rect 294414 70252 294420 70304
rect 294472 70292 294478 70304
rect 295978 70292 295984 70304
rect 294472 70264 295984 70292
rect 294472 70252 294478 70264
rect 295978 70252 295984 70264
rect 296036 70252 296042 70304
rect 296073 70295 296131 70301
rect 296073 70261 296085 70295
rect 296119 70292 296131 70295
rect 325786 70292 325792 70304
rect 296119 70264 325792 70292
rect 296119 70261 296131 70264
rect 296073 70255 296131 70261
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 325786 70252 325792 70264
rect 325844 70252 325850 70304
rect 338022 70252 338028 70304
rect 338080 70292 338086 70304
rect 353754 70292 353760 70304
rect 338080 70264 353760 70292
rect 338080 70252 338086 70264
rect 353754 70252 353760 70264
rect 353812 70252 353818 70304
<<<<<<< HEAD
rect 378226 70252 378232 70304
rect 378284 70292 378290 70304
rect 388441 70295 388499 70301
rect 378284 70264 383976 70292
rect 378284 70252 378290 70264
=======
rect 375374 70252 375380 70304
rect 375432 70292 375438 70304
rect 447134 70292 447140 70304
rect 375432 70264 447140 70292
rect 375432 70252 375438 70264
rect 447134 70252 447140 70264
rect 447192 70252 447198 70304
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 34422 70184 34428 70236
rect 34480 70224 34486 70236
rect 59449 70227 59507 70233
rect 59449 70224 59461 70227
rect 34480 70196 59461 70224
rect 34480 70184 34486 70196
rect 59449 70193 59461 70196
rect 59495 70193 59507 70227
rect 59449 70187 59507 70193
rect 59541 70227 59599 70233
rect 59541 70193 59553 70227
rect 59587 70224 59599 70227
rect 64874 70224 64880 70236
rect 59587 70196 64880 70224
rect 59587 70193 59599 70196
rect 59541 70187 59599 70193
rect 64874 70184 64880 70196
rect 64932 70184 64938 70236
rect 84378 70224 84384 70236
rect 74506 70196 84384 70224
rect 50338 70116 50344 70168
rect 50396 70156 50402 70168
rect 74506 70156 74534 70196
rect 84378 70184 84384 70196
rect 84436 70184 84442 70236
rect 119338 70184 119344 70236
rect 119396 70224 119402 70236
rect 127618 70224 127624 70236
rect 119396 70196 127624 70224
rect 119396 70184 119402 70196
rect 127618 70184 127624 70196
rect 127676 70184 127682 70236
rect 144822 70184 144828 70236
rect 144880 70224 144886 70236
rect 226702 70224 226708 70236
rect 144880 70196 226708 70224
rect 144880 70184 144886 70196
rect 226702 70184 226708 70196
rect 226760 70184 226766 70236
rect 291654 70184 291660 70236
rect 291712 70224 291718 70236
<<<<<<< HEAD
rect 300857 70227 300915 70233
rect 300857 70224 300869 70227
rect 291712 70196 300869 70224
rect 291712 70184 291718 70196
rect 300857 70193 300869 70196
rect 300903 70193 300915 70227
rect 300857 70187 300915 70193
rect 301501 70227 301559 70233
rect 301501 70193 301513 70227
rect 301547 70224 301559 70227
rect 345382 70224 345388 70236
rect 301547 70196 345388 70224
rect 301547 70193 301559 70196
rect 301501 70187 301559 70193
rect 345382 70184 345388 70196
rect 345440 70184 345446 70236
rect 380986 70184 380992 70236
rect 381044 70224 381050 70236
rect 383841 70227 383899 70233
rect 383841 70224 383853 70227
rect 381044 70196 383853 70224
rect 381044 70184 381050 70196
rect 383841 70193 383853 70196
rect 383887 70193 383899 70227
rect 383948 70224 383976 70264
rect 388441 70261 388453 70295
rect 388487 70292 388499 70295
rect 454034 70292 454040 70304
rect 388487 70264 454040 70292
rect 388487 70261 388499 70264
rect 388441 70255 388499 70261
rect 454034 70252 454040 70264
rect 454092 70252 454098 70304
rect 460934 70224 460940 70236
rect 383948 70196 460940 70224
rect 383841 70187 383899 70193
rect 460934 70184 460940 70196
rect 460992 70184 460998 70236
=======
rect 301501 70227 301559 70233
rect 301501 70224 301513 70227
rect 291712 70196 301513 70224
rect 291712 70184 291718 70196
rect 301501 70193 301513 70196
rect 301547 70193 301559 70227
rect 301501 70187 301559 70193
rect 301593 70227 301651 70233
rect 301593 70193 301605 70227
rect 301639 70224 301651 70227
rect 345382 70224 345388 70236
rect 301639 70196 345388 70224
rect 301639 70193 301651 70196
rect 301593 70187 301651 70193
rect 345382 70184 345388 70196
rect 345440 70184 345446 70236
rect 379606 70184 379612 70236
rect 379664 70224 379670 70236
rect 388533 70227 388591 70233
rect 388533 70224 388545 70227
rect 379664 70196 388545 70224
rect 379664 70184 379670 70196
rect 388533 70193 388545 70196
rect 388579 70193 388591 70227
rect 388533 70187 388591 70193
rect 388625 70227 388683 70233
rect 388625 70193 388637 70227
rect 388671 70224 388683 70227
rect 454034 70224 454040 70236
rect 388671 70196 454040 70224
rect 388671 70193 388683 70196
rect 388625 70187 388683 70193
rect 454034 70184 454040 70196
rect 454092 70184 454098 70236
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 50396 70128 74534 70156
rect 50396 70116 50402 70128
rect 80882 70116 80888 70168
rect 80940 70156 80946 70168
rect 88337 70159 88395 70165
rect 88337 70156 88349 70159
rect 80940 70128 88349 70156
rect 80940 70116 80946 70128
rect 88337 70125 88349 70128
rect 88383 70125 88395 70159
rect 95510 70156 95516 70168
rect 88337 70119 88395 70125
rect 93826 70128 95516 70156
rect 27522 70048 27528 70100
rect 27580 70088 27586 70100
rect 59541 70091 59599 70097
rect 59541 70088 59553 70091
rect 27580 70060 59553 70088
rect 27580 70048 27586 70060
rect 59541 70057 59553 70060
rect 59587 70057 59599 70091
rect 59541 70051 59599 70057
rect 68278 70048 68284 70100
rect 68336 70088 68342 70100
rect 93826 70088 93854 70128
rect 95510 70116 95516 70128
rect 95568 70116 95574 70168
rect 106734 70116 106740 70168
rect 106792 70156 106798 70168
rect 122834 70156 122840 70168
rect 106792 70128 122840 70156
rect 106792 70116 106798 70128
rect 122834 70116 122840 70128
rect 122892 70116 122898 70168
rect 137922 70116 137928 70168
rect 137980 70156 137986 70168
rect 225322 70156 225328 70168
rect 137980 70128 225328 70156
rect 137980 70116 137986 70128
rect 225322 70116 225328 70128
rect 225380 70116 225386 70168
rect 231118 70116 231124 70168
rect 231176 70156 231182 70168
rect 239950 70156 239956 70168
rect 231176 70128 239956 70156
rect 231176 70116 231182 70128
rect 239950 70116 239956 70128
rect 240008 70116 240014 70168
<<<<<<< HEAD
rect 281442 70116 281448 70168
rect 281500 70156 281506 70168
rect 342346 70156 342352 70168
rect 281500 70128 342352 70156
rect 281500 70116 281506 70128
rect 342346 70116 342352 70128
rect 342404 70116 342410 70168
rect 379606 70116 379612 70168
rect 379664 70156 379670 70168
rect 467834 70156 467840 70168
rect 379664 70128 467840 70156
rect 379664 70116 379670 70128
rect 467834 70116 467840 70128
rect 467892 70116 467898 70168
=======
rect 250346 70156 250352 70168
rect 248386 70128 250352 70156
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 68336 70060 93854 70088
rect 68336 70048 68342 70060
rect 103422 70048 103428 70100
rect 103480 70088 103486 70100
rect 103480 70048 103514 70088
rect 107470 70048 107476 70100
rect 107528 70088 107534 70100
rect 125594 70088 125600 70100
rect 107528 70060 125600 70088
rect 107528 70048 107534 70060
rect 125594 70048 125600 70060
rect 125652 70048 125658 70100
rect 163958 70048 163964 70100
rect 164016 70088 164022 70100
<<<<<<< HEAD
rect 250346 70088 250352 70100
rect 164016 70060 250352 70088
rect 164016 70048 164022 70060
rect 250346 70048 250352 70060
rect 250404 70048 250410 70100
=======
rect 248386 70088 248414 70128
rect 250346 70116 250352 70128
rect 250404 70116 250410 70168
rect 281442 70116 281448 70168
rect 281500 70156 281506 70168
rect 342346 70156 342352 70168
rect 281500 70128 342352 70156
rect 281500 70116 281506 70128
rect 342346 70116 342352 70128
rect 342404 70116 342410 70168
rect 378226 70116 378232 70168
rect 378284 70156 378290 70168
rect 460934 70156 460940 70168
rect 378284 70128 460940 70156
rect 378284 70116 378290 70128
rect 460934 70116 460940 70128
rect 460992 70116 460998 70168
rect 164016 70060 248414 70088
rect 164016 70048 164022 70060
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 295794 70048 295800 70100
rect 295852 70088 295858 70100
rect 410518 70088 410524 70100
rect 295852 70060 410524 70088
rect 295852 70048 295858 70060
rect 410518 70048 410524 70060
rect 410576 70048 410582 70100
rect 51718 69980 51724 70032
rect 51776 70020 51782 70032
rect 92014 70020 92020 70032
rect 51776 69992 92020 70020
rect 51776 69980 51782 69992
rect 92014 69980 92020 69992
rect 92072 69980 92078 70032
rect 103486 70020 103514 70048
rect 124858 70020 124864 70032
rect 103486 69992 124864 70020
rect 124858 69980 124864 69992
rect 124916 69980 124922 70032
rect 135162 69980 135168 70032
rect 135220 70020 135226 70032
rect 224678 70020 224684 70032
rect 135220 69992 224684 70020
rect 135220 69980 135226 69992
rect 224678 69980 224684 69992
rect 224736 69980 224742 70032
rect 234522 69980 234528 70032
rect 234580 70020 234586 70032
rect 244182 70020 244188 70032
rect 234580 69992 244188 70020
rect 234580 69980 234586 69992
rect 244182 69980 244188 69992
rect 244240 69980 244246 70032
rect 295150 69980 295156 70032
rect 295208 70020 295214 70032
rect 418798 70020 418804 70032
rect 295208 69992 418804 70020
rect 295208 69980 295214 69992
rect 418798 69980 418804 69992
rect 418856 69980 418862 70032
rect 17862 69912 17868 69964
rect 17920 69952 17926 69964
rect 63494 69952 63500 69964
rect 17920 69924 63500 69952
rect 17920 69912 17926 69924
rect 63494 69912 63500 69924
rect 63552 69912 63558 69964
rect 88337 69955 88395 69961
rect 88337 69921 88349 69955
rect 88383 69952 88395 69955
rect 107562 69952 107568 69964
rect 88383 69924 107568 69952
rect 88383 69921 88395 69924
rect 88337 69915 88395 69921
rect 107562 69912 107568 69924
rect 107620 69912 107626 69964
rect 114462 69912 114468 69964
rect 114520 69952 114526 69964
rect 126974 69952 126980 69964
rect 114520 69924 126980 69952
rect 114520 69912 114526 69924
rect 126974 69912 126980 69924
rect 127032 69912 127038 69964
<<<<<<< HEAD
rect 204901 69955 204959 69961
rect 204901 69921 204913 69955
rect 204947 69952 204959 69955
rect 353938 69952 353944 69964
rect 204947 69924 353944 69952
rect 204947 69921 204959 69924
rect 204901 69915 204959 69921
rect 353938 69912 353944 69924
rect 353996 69912 354002 69964
rect 383841 69955 383899 69961
rect 383841 69921 383853 69955
rect 383887 69952 383899 69955
rect 474734 69952 474740 69964
rect 383887 69924 474740 69952
rect 383887 69921 383899 69924
rect 383841 69915 383899 69921
rect 474734 69912 474740 69924
rect 474792 69912 474798 69964
=======
rect 204809 69955 204867 69961
rect 204809 69921 204821 69955
rect 204855 69952 204867 69955
rect 353938 69952 353944 69964
rect 204855 69924 353944 69952
rect 204855 69921 204867 69924
rect 204809 69915 204867 69921
rect 353938 69912 353944 69924
rect 353996 69912 354002 69964
rect 380986 69912 380992 69964
rect 381044 69952 381050 69964
rect 388533 69955 388591 69961
rect 381044 69924 388484 69952
rect 381044 69912 381050 69924
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 7558 69844 7564 69896
rect 7616 69884 7622 69896
rect 60274 69884 60280 69896
rect 7616 69856 60280 69884
rect 7616 69844 7622 69856
rect 60274 69844 60280 69856
rect 60332 69844 60338 69896
rect 65518 69844 65524 69896
rect 65576 69884 65582 69896
rect 92474 69884 92480 69896
rect 65576 69856 92480 69884
rect 65576 69844 65582 69856
rect 92474 69844 92480 69856
rect 92532 69844 92538 69896
rect 93118 69844 93124 69896
rect 93176 69884 93182 69896
rect 94130 69884 94136 69896
rect 93176 69856 94136 69884
rect 93176 69844 93182 69856
rect 94130 69844 94136 69856
rect 94188 69844 94194 69896
rect 103238 69844 103244 69896
rect 103296 69884 103302 69896
rect 104158 69884 104164 69896
rect 103296 69856 104164 69884
rect 103296 69844 103302 69856
rect 104158 69844 104164 69856
rect 104216 69844 104222 69896
rect 108301 69887 108359 69893
rect 108301 69853 108313 69887
rect 108347 69884 108359 69887
rect 124122 69884 124128 69896
rect 108347 69856 124128 69884
rect 108347 69853 108359 69856
rect 108301 69847 108359 69853
rect 124122 69844 124128 69856
rect 124180 69844 124186 69896
<<<<<<< HEAD
rect 131022 69844 131028 69896
rect 131080 69884 131086 69896
rect 223942 69884 223948 69896
rect 131080 69856 223948 69884
rect 131080 69844 131086 69856
rect 223942 69844 223948 69856
rect 224000 69844 224006 69896
rect 228358 69844 228364 69896
rect 228416 69884 228422 69896
rect 230198 69884 230204 69896
rect 228416 69856 230204 69884
rect 228416 69844 228422 69856
rect 230198 69844 230204 69856
rect 230256 69844 230262 69896
rect 230477 69887 230535 69893
rect 230477 69853 230489 69887
rect 230523 69884 230535 69887
rect 242802 69884 242808 69896
rect 230523 69856 242808 69884
rect 230523 69853 230535 69856
rect 230477 69847 230535 69853
rect 242802 69844 242808 69856
rect 242860 69844 242866 69896
rect 250438 69844 250444 69896
rect 250496 69884 250502 69896
rect 264974 69884 264980 69896
rect 250496 69856 264980 69884
rect 250496 69844 250502 69856
rect 264974 69844 264980 69856
rect 265032 69844 265038 69896
rect 300857 69887 300915 69893
rect 300857 69853 300869 69887
rect 300903 69884 300915 69887
rect 472618 69884 472624 69896
rect 300903 69856 472624 69884
rect 300903 69853 300915 69856
rect 300857 69847 300915 69853
rect 472618 69844 472624 69856
rect 472676 69844 472682 69896
=======
rect 129642 69844 129648 69896
rect 129700 69884 129706 69896
rect 134610 69884 134616 69896
rect 129700 69856 134616 69884
rect 129700 69844 129706 69856
rect 134610 69844 134616 69856
rect 134668 69844 134674 69896
rect 213457 69887 213515 69893
rect 200086 69856 209774 69884
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 18598 69776 18604 69828
rect 18656 69816 18662 69828
rect 107654 69816 107660 69828
rect 18656 69788 107660 69816
rect 18656 69776 18662 69788
rect 107654 69776 107660 69788
rect 107712 69776 107718 69828
rect 111702 69776 111708 69828
rect 111760 69816 111766 69828
rect 126238 69816 126244 69828
rect 111760 69788 126244 69816
rect 111760 69776 111766 69788
rect 126238 69776 126244 69788
rect 126296 69776 126302 69828
<<<<<<< HEAD
rect 129642 69776 129648 69828
rect 129700 69816 129706 69828
rect 134610 69816 134616 69828
rect 129700 69788 134616 69816
rect 129700 69776 129706 69788
rect 134610 69776 134616 69788
rect 134668 69776 134674 69828
rect 154206 69776 154212 69828
rect 154264 69816 154270 69828
rect 204990 69816 204996 69828
rect 154264 69788 204996 69816
rect 154264 69776 154270 69788
rect 204990 69776 204996 69788
rect 205048 69776 205054 69828
rect 208578 69776 208584 69828
rect 208636 69816 208642 69828
rect 413278 69816 413284 69828
rect 208636 69788 413284 69816
rect 208636 69776 208642 69788
rect 413278 69776 413284 69788
rect 413336 69776 413342 69828
=======
rect 131022 69776 131028 69828
rect 131080 69816 131086 69828
rect 200086 69816 200114 69856
rect 131080 69788 200114 69816
rect 209746 69816 209774 69856
rect 213457 69853 213469 69887
rect 213503 69884 213515 69887
rect 371786 69884 371792 69896
rect 213503 69856 371792 69884
rect 213503 69853 213515 69856
rect 213457 69847 213515 69853
rect 371786 69844 371792 69856
rect 371844 69844 371850 69896
rect 388456 69884 388484 69924
rect 388533 69921 388545 69955
rect 388579 69952 388591 69955
rect 467834 69952 467840 69964
rect 388579 69924 467840 69952
rect 388579 69921 388591 69924
rect 388533 69915 388591 69921
rect 467834 69912 467840 69924
rect 467892 69912 467898 69964
rect 474734 69884 474740 69896
rect 388456 69856 474740 69884
rect 474734 69844 474740 69856
rect 474792 69844 474798 69896
rect 223942 69816 223948 69828
rect 209746 69788 223948 69816
rect 131080 69776 131086 69788
rect 223942 69776 223948 69788
rect 224000 69776 224006 69828
rect 228358 69776 228364 69828
rect 228416 69816 228422 69828
rect 230198 69816 230204 69828
rect 228416 69788 230204 69816
rect 228416 69776 228422 69788
rect 230198 69776 230204 69788
rect 230256 69776 230262 69828
rect 233789 69819 233847 69825
rect 233789 69785 233801 69819
rect 233835 69816 233847 69819
rect 242802 69816 242808 69828
rect 233835 69788 242808 69816
rect 233835 69785 233847 69788
rect 233789 69779 233847 69785
rect 242802 69776 242808 69788
rect 242860 69776 242866 69828
rect 250438 69776 250444 69828
rect 250496 69816 250502 69828
rect 264974 69816 264980 69828
rect 250496 69788 264980 69816
rect 250496 69776 250502 69788
rect 264974 69776 264980 69788
rect 265032 69776 265038 69828
rect 287698 69776 287704 69828
rect 287756 69816 287762 69828
rect 296073 69819 296131 69825
rect 296073 69816 296085 69819
rect 287756 69788 296085 69816
rect 287756 69776 287762 69788
rect 296073 69785 296085 69788
rect 296119 69785 296131 69819
rect 296073 69779 296131 69785
rect 301501 69819 301559 69825
rect 301501 69785 301513 69819
rect 301547 69816 301559 69819
rect 472618 69816 472624 69828
rect 301547 69788 472624 69816
rect 301547 69785 301559 69788
rect 301501 69779 301559 69785
rect 472618 69776 472624 69788
rect 472676 69776 472682 69828
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 21358 69708 21364 69760
rect 21416 69748 21422 69760
rect 130470 69748 130476 69760
rect 21416 69720 130476 69748
rect 21416 69708 21422 69720
rect 130470 69708 130476 69720
rect 130528 69708 130534 69760
<<<<<<< HEAD
rect 209961 69751 210019 69757
rect 209961 69717 209973 69751
rect 210007 69748 210019 69751
rect 411898 69748 411904 69760
rect 210007 69720 411904 69748
rect 210007 69717 210019 69720
rect 209961 69711 210019 69717
rect 411898 69708 411904 69720
rect 411956 69708 411962 69760
=======
rect 154206 69708 154212 69760
rect 154264 69748 154270 69760
rect 204898 69748 204904 69760
rect 154264 69720 204904 69748
rect 154264 69708 154270 69720
rect 204898 69708 204904 69720
rect 204956 69708 204962 69760
rect 208578 69708 208584 69760
rect 208636 69748 208642 69760
rect 413278 69748 413284 69760
rect 208636 69720 413284 69748
rect 208636 69708 208642 69720
rect 413278 69708 413284 69720
rect 413336 69708 413342 69760
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 11698 69640 11704 69692
rect 11756 69680 11762 69692
rect 133230 69680 133236 69692
rect 11756 69652 133236 69680
rect 11756 69640 11762 69652
rect 133230 69640 133236 69652
rect 133288 69640 133294 69692
rect 193306 69640 193312 69692
rect 193364 69680 193370 69692
<<<<<<< HEAD
rect 204901 69683 204959 69689
rect 204901 69680 204913 69683
rect 193364 69652 204913 69680
rect 193364 69640 193370 69652
rect 204901 69649 204913 69652
rect 204947 69649 204959 69683
rect 204901 69643 204959 69649
rect 205082 69640 205088 69692
rect 205140 69680 205146 69692
rect 371786 69680 371792 69692
rect 205140 69652 371792 69680
rect 205140 69640 205146 69652
rect 371786 69640 371792 69652
rect 371844 69640 371850 69692
rect 376754 69640 376760 69692
rect 376812 69680 376818 69692
rect 388441 69683 388499 69689
rect 388441 69680 388453 69683
rect 376812 69652 388453 69680
rect 376812 69640 376818 69652
rect 388441 69649 388453 69652
rect 388487 69649 388499 69683
rect 388441 69643 388499 69649
=======
rect 204809 69683 204867 69689
rect 204809 69680 204821 69683
rect 193364 69652 204821 69680
rect 193364 69640 193370 69652
rect 204809 69649 204821 69652
rect 204855 69649 204867 69683
rect 204809 69643 204867 69649
rect 205082 69640 205088 69692
rect 205140 69680 205146 69692
rect 213457 69683 213515 69689
rect 213457 69680 213469 69683
rect 205140 69652 213469 69680
rect 205140 69640 205146 69652
rect 213457 69649 213469 69652
rect 213503 69649 213515 69683
rect 213457 69643 213515 69649
rect 214561 69683 214619 69689
rect 214561 69649 214573 69683
rect 214607 69680 214619 69683
rect 411898 69680 411904 69692
rect 214607 69652 411904 69680
rect 214607 69649 214619 69652
rect 214561 69643 214619 69649
rect 411898 69640 411904 69652
rect 411956 69640 411962 69692
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 59449 69615 59507 69621
rect 59449 69581 59461 69615
rect 59495 69612 59507 69615
rect 66254 69612 66260 69624
rect 59495 69584 66260 69612
rect 59495 69581 59507 69584
rect 59449 69575 59507 69581
rect 66254 69572 66260 69584
rect 66312 69572 66318 69624
rect 81618 69572 81624 69624
rect 81676 69612 81682 69624
rect 86218 69612 86224 69624
rect 81676 69584 86224 69612
rect 81676 69572 81682 69584
rect 86218 69572 86224 69584
rect 86276 69572 86282 69624
rect 100662 69572 100668 69624
rect 100720 69612 100726 69624
rect 108301 69615 108359 69621
rect 108301 69612 108313 69615
rect 100720 69584 108313 69612
rect 100720 69572 100726 69584
rect 108301 69581 108313 69584
rect 108347 69581 108359 69615
rect 108301 69575 108359 69581
rect 155862 69572 155868 69624
rect 155920 69612 155926 69624
rect 155920 69584 224356 69612
rect 155920 69572 155926 69584
rect 65886 69504 65892 69556
rect 65944 69544 65950 69556
rect 66898 69544 66904 69556
rect 65944 69516 66904 69544
rect 65944 69504 65950 69516
rect 66898 69504 66904 69516
rect 66956 69504 66962 69556
rect 157702 69504 157708 69556
rect 157760 69544 157766 69556
rect 224218 69544 224224 69556
rect 157760 69516 224224 69544
rect 157760 69504 157766 69516
rect 224218 69504 224224 69516
rect 224276 69504 224282 69556
rect 224328 69544 224356 69584
rect 227622 69572 227628 69624
rect 227680 69612 227686 69624
<<<<<<< HEAD
rect 230477 69615 230535 69621
rect 230477 69612 230489 69615
rect 227680 69584 230489 69612
rect 227680 69572 227686 69584
rect 230477 69581 230489 69584
rect 230523 69581 230535 69615
rect 230477 69575 230535 69581
=======
rect 233789 69615 233847 69621
rect 233789 69612 233801 69615
rect 227680 69584 233801 69612
rect 227680 69572 227686 69584
rect 233789 69581 233801 69584
rect 233835 69581 233847 69615
rect 233789 69575 233847 69581
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 247678 69572 247684 69624
rect 247736 69612 247742 69624
rect 248966 69612 248972 69624
rect 247736 69584 248972 69612
rect 247736 69572 247742 69584
rect 248966 69572 248972 69584
rect 249024 69572 249030 69624
<<<<<<< HEAD
rect 272150 69572 272156 69624
rect 272208 69612 272214 69624
rect 274358 69612 274364 69624
rect 272208 69584 274364 69612
rect 272208 69572 272214 69584
rect 274358 69572 274364 69584
rect 274416 69572 274422 69624
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 293770 69572 293776 69624
rect 293828 69612 293834 69624
rect 310146 69612 310152 69624
rect 293828 69584 310152 69612
rect 293828 69572 293834 69584
rect 310146 69572 310152 69584
rect 310204 69572 310210 69624
rect 313182 69572 313188 69624
rect 313240 69612 313246 69624
rect 348878 69612 348884 69624
rect 313240 69584 348884 69612
rect 313240 69572 313246 69584
rect 348878 69572 348884 69584
rect 348936 69572 348942 69624
<<<<<<< HEAD
rect 373994 69572 374000 69624
rect 374052 69612 374058 69624
rect 440234 69612 440240 69624
rect 374052 69584 440240 69612
rect 374052 69572 374058 69584
rect 440234 69572 440240 69584
rect 440292 69572 440298 69624
=======
rect 372614 69572 372620 69624
rect 372672 69612 372678 69624
rect 431954 69612 431960 69624
rect 372672 69584 431960 69612
rect 372672 69572 372678 69584
rect 431954 69572 431960 69584
rect 432012 69572 432018 69624
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 228818 69544 228824 69556
rect 224328 69516 228824 69544
rect 228818 69504 228824 69516
rect 228876 69504 228882 69556
rect 291838 69504 291844 69556
rect 291896 69544 291902 69556
rect 323026 69544 323032 69556
rect 291896 69516 323032 69544
rect 291896 69504 291902 69516
rect 323026 69504 323032 69516
rect 323084 69504 323090 69556
rect 324222 69504 324228 69556
rect 324280 69544 324286 69556
rect 350626 69544 350632 69556
rect 324280 69516 350632 69544
rect 324280 69504 324286 69516
rect 350626 69504 350632 69516
rect 350684 69504 350690 69556
<<<<<<< HEAD
rect 372614 69504 372620 69556
rect 372672 69544 372678 69556
rect 431954 69544 431960 69556
rect 372672 69516 431960 69544
rect 372672 69504 372678 69516
rect 431954 69504 431960 69516
rect 432012 69504 432018 69556
=======
rect 371878 69504 371884 69556
rect 371936 69544 371942 69556
rect 429194 69544 429200 69556
rect 371936 69516 429200 69544
rect 371936 69504 371942 69516
rect 429194 69504 429200 69516
rect 429252 69504 429258 69556
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 164694 69436 164700 69488
rect 164752 69476 164758 69488
rect 226978 69476 226984 69488
rect 164752 69448 226984 69476
rect 164752 69436 164758 69448
rect 226978 69436 226984 69448
rect 227036 69436 227042 69488
<<<<<<< HEAD
=======
rect 272150 69436 272156 69488
rect 272208 69476 272214 69488
rect 274358 69476 274364 69488
rect 272208 69448 274364 69476
rect 272208 69436 272214 69448
rect 274358 69436 274364 69448
rect 274416 69436 274422 69488
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 289078 69436 289084 69488
rect 289136 69476 289142 69488
rect 320266 69476 320272 69488
rect 289136 69448 320272 69476
rect 289136 69436 289142 69448
rect 320266 69436 320272 69448
rect 320324 69436 320330 69488
rect 342162 69436 342168 69488
rect 342220 69476 342226 69488
rect 354398 69476 354404 69488
rect 342220 69448 354404 69476
rect 342220 69436 342226 69448
rect 354398 69436 354404 69448
rect 354456 69436 354462 69488
<<<<<<< HEAD
rect 371878 69436 371884 69488
rect 371936 69476 371942 69488
rect 429194 69476 429200 69488
rect 371936 69448 429200 69476
rect 371936 69436 371942 69448
rect 429194 69436 429200 69448
rect 429252 69436 429258 69488
=======
rect 370498 69436 370504 69488
rect 370556 69476 370562 69488
rect 422294 69476 422300 69488
rect 370556 69448 422300 69476
rect 370556 69436 370562 69448
rect 422294 69436 422300 69448
rect 422352 69436 422358 69488
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 126882 69368 126888 69420
rect 126940 69408 126946 69420
rect 133874 69408 133880 69420
rect 126940 69380 133880 69408
rect 126940 69368 126946 69380
rect 133874 69368 133880 69380
rect 133932 69368 133938 69420
rect 154850 69368 154856 69420
rect 154908 69408 154914 69420
rect 206278 69408 206284 69420
rect 154908 69380 206284 69408
rect 154908 69368 154914 69380
rect 206278 69368 206284 69380
rect 206336 69368 206342 69420
rect 209682 69368 209688 69420
rect 209740 69408 209746 69420
rect 239306 69408 239312 69420
rect 209740 69380 239312 69408
rect 209740 69368 209746 69380
rect 239306 69368 239312 69380
rect 239364 69368 239370 69420
rect 293034 69368 293040 69420
rect 293092 69408 293098 69420
rect 310330 69408 310336 69420
rect 293092 69380 310336 69408
rect 293092 69368 293098 69380
rect 310330 69368 310336 69380
rect 310388 69368 310394 69420
<<<<<<< HEAD
rect 370498 69368 370504 69420
rect 370556 69408 370562 69420
rect 422294 69408 422300 69420
rect 370556 69380 422300 69408
rect 370556 69368 370562 69380
rect 422294 69368 422300 69380
rect 422352 69368 422358 69420
=======
rect 367738 69368 367744 69420
rect 367796 69408 367802 69420
rect 407114 69408 407120 69420
rect 367796 69380 407120 69408
rect 367796 69368 367802 69380
rect 407114 69368 407120 69380
rect 407172 69368 407178 69420
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 156322 69300 156328 69352
rect 156380 69340 156386 69352
rect 204898 69340 204904 69352
rect 156380 69312 204904 69340
rect 156380 69300 156386 69312
rect 204898 69300 204904 69312
rect 204956 69300 204962 69352
rect 207198 69300 207204 69352
rect 207256 69340 207262 69352
rect 224310 69340 224316 69352
rect 207256 69312 224316 69340
rect 207256 69300 207262 69312
rect 224310 69300 224316 69312
rect 224368 69300 224374 69352
rect 290274 69300 290280 69352
rect 290332 69340 290338 69352
rect 292390 69340 292396 69352
rect 290332 69312 292396 69340
rect 290332 69300 290338 69312
rect 292390 69300 292396 69312
rect 292448 69300 292454 69352
rect 295242 69300 295248 69352
rect 295300 69340 295306 69352
<<<<<<< HEAD
rect 301501 69343 301559 69349
rect 301501 69340 301513 69343
rect 295300 69312 301513 69340
rect 295300 69300 295306 69312
rect 301501 69309 301513 69312
rect 301547 69309 301559 69343
rect 301501 69303 301559 69309
rect 367738 69300 367744 69352
rect 367796 69340 367802 69352
rect 407114 69340 407120 69352
rect 367796 69312 407120 69340
rect 367796 69300 367802 69312
rect 407114 69300 407120 69312
rect 407172 69300 407178 69352
=======
rect 301593 69343 301651 69349
rect 301593 69340 301605 69343
rect 295300 69312 301605 69340
rect 295300 69300 295306 69312
rect 301593 69309 301605 69312
rect 301639 69309 301651 69343
rect 301593 69303 301651 69309
rect 376754 69300 376760 69352
rect 376812 69340 376818 69352
rect 388625 69343 388683 69349
rect 388625 69340 388637 69343
rect 376812 69312 388637 69340
rect 376812 69300 376818 69312
rect 388625 69309 388637 69312
rect 388671 69309 388683 69343
rect 414658 69340 414664 69352
rect 388625 69303 388683 69309
rect 393286 69312 414664 69340
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 111794 69232 111800 69284
rect 111852 69272 111858 69284
rect 114370 69272 114376 69284
rect 111852 69244 114376 69272
rect 111852 69232 111858 69244
rect 114370 69232 114376 69244
rect 114428 69232 114434 69284
rect 163222 69232 163228 69284
rect 163280 69272 163286 69284
rect 209130 69272 209136 69284
rect 163280 69244 209136 69272
rect 163280 69232 163286 69244
rect 209130 69232 209136 69244
rect 209188 69232 209194 69284
<<<<<<< HEAD
=======
rect 209961 69275 210019 69281
rect 209961 69241 209973 69275
rect 210007 69272 210019 69275
rect 214561 69275 214619 69281
rect 214561 69272 214573 69275
rect 210007 69244 214573 69272
rect 210007 69241 210019 69244
rect 209961 69235 210019 69241
rect 214561 69241 214573 69244
rect 214607 69241 214619 69275
rect 214561 69235 214619 69241
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 222838 69232 222844 69284
rect 222896 69272 222902 69284
rect 233234 69272 233240 69284
rect 222896 69244 233240 69272
rect 222896 69232 222902 69244
rect 233234 69232 233240 69244
rect 233292 69232 233298 69284
<<<<<<< HEAD
rect 294414 69232 294420 69284
rect 294472 69272 294478 69284
rect 295886 69272 295892 69284
rect 294472 69244 295892 69272
rect 294472 69232 294478 69244
rect 295886 69232 295892 69244
rect 295944 69232 295950 69284
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 309870 69232 309876 69284
rect 309928 69272 309934 69284
rect 319530 69272 319536 69284
rect 309928 69244 319536 69272
rect 309928 69232 309934 69244
rect 319530 69232 319536 69244
rect 319588 69232 319594 69284
rect 383746 69232 383752 69284
rect 383804 69272 383810 69284
<<<<<<< HEAD
rect 414658 69272 414664 69284
rect 383804 69244 414664 69272
rect 383804 69232 383810 69244
rect 414658 69232 414664 69244
rect 414716 69232 414722 69284
=======
rect 393286 69272 393314 69312
rect 414658 69300 414664 69312
rect 414716 69300 414722 69352
rect 383804 69244 393314 69272
rect 383804 69232 383810 69244
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 78122 69164 78128 69216
rect 78180 69204 78186 69216
rect 83458 69204 83464 69216
rect 78180 69176 83464 69204
rect 78180 69164 78186 69176
rect 83458 69164 83464 69176
rect 83516 69164 83522 69216
rect 197998 69164 198004 69216
rect 198056 69204 198062 69216
rect 236454 69204 236460 69216
rect 198056 69176 236460 69204
rect 198056 69164 198062 69176
rect 236454 69164 236460 69176
rect 236512 69164 236518 69216
rect 57238 69096 57244 69148
rect 57296 69136 57302 69148
rect 61378 69136 61384 69148
rect 57296 69108 61384 69136
rect 57296 69096 57302 69108
rect 61378 69096 61384 69108
rect 61436 69096 61442 69148
rect 72418 69096 72424 69148
rect 72476 69136 72482 69148
rect 73246 69136 73252 69148
rect 72476 69108 73252 69136
rect 72476 69096 72482 69108
rect 73246 69096 73252 69108
rect 73304 69096 73310 69148
rect 74626 69096 74632 69148
rect 74684 69136 74690 69148
rect 75730 69136 75736 69148
rect 74684 69108 75736 69136
rect 74684 69096 74690 69108
rect 75730 69096 75736 69108
rect 75788 69096 75794 69148
rect 76006 69096 76012 69148
rect 76064 69136 76070 69148
rect 77110 69136 77116 69148
rect 76064 69108 77116 69136
rect 76064 69096 76070 69108
rect 77110 69096 77116 69108
rect 77168 69096 77174 69148
rect 78858 69096 78864 69148
rect 78916 69136 78922 69148
rect 79962 69136 79968 69148
rect 78916 69108 79968 69136
rect 78916 69096 78922 69108
rect 79962 69096 79968 69108
rect 80020 69096 80026 69148
rect 94498 69096 94504 69148
rect 94556 69136 94562 69148
rect 100386 69136 100392 69148
rect 94556 69108 100392 69136
rect 94556 69096 94562 69108
rect 100386 69096 100392 69108
rect 100444 69096 100450 69148
rect 173066 69096 173072 69148
rect 173124 69136 173130 69148
rect 173802 69136 173808 69148
rect 173124 69108 173808 69136
rect 173124 69096 173130 69108
rect 173802 69096 173808 69108
rect 173860 69096 173866 69148
rect 186314 69096 186320 69148
rect 186372 69136 186378 69148
rect 187602 69136 187608 69148
rect 186372 69108 187608 69136
rect 186372 69096 186378 69108
rect 187602 69096 187608 69108
rect 187660 69096 187666 69148
rect 187694 69096 187700 69148
rect 187752 69136 187758 69148
rect 188890 69136 188896 69148
rect 187752 69108 188896 69136
rect 187752 69096 187758 69108
rect 188890 69096 188896 69108
rect 188948 69096 188954 69148
rect 189074 69096 189080 69148
rect 189132 69136 189138 69148
rect 190270 69136 190276 69148
rect 189132 69108 190276 69136
rect 189132 69096 189138 69108
rect 190270 69096 190276 69108
rect 190328 69096 190334 69148
rect 190454 69096 190460 69148
rect 190512 69136 190518 69148
rect 191650 69136 191656 69148
rect 190512 69108 191656 69136
rect 190512 69096 190518 69108
rect 191650 69096 191656 69108
rect 191708 69096 191714 69148
rect 194686 69096 194692 69148
rect 194744 69136 194750 69148
rect 195882 69136 195888 69148
rect 194744 69108 195888 69136
rect 194744 69096 194750 69108
rect 195882 69096 195888 69108
rect 195940 69096 195946 69148
rect 196066 69096 196072 69148
rect 196124 69136 196130 69148
rect 197170 69136 197176 69148
rect 196124 69108 197176 69136
rect 196124 69096 196130 69108
rect 197170 69096 197176 69108
rect 197228 69096 197234 69148
rect 198826 69096 198832 69148
rect 198884 69136 198890 69148
rect 199930 69136 199936 69148
rect 198884 69108 199936 69136
rect 198884 69096 198890 69108
rect 199930 69096 199936 69108
rect 199988 69096 199994 69148
rect 203702 69096 203708 69148
rect 203760 69136 203766 69148
rect 203760 69108 206784 69136
rect 203760 69096 203766 69108
rect 58618 69028 58624 69080
rect 58676 69068 58682 69080
rect 60642 69068 60648 69080
rect 58676 69040 60648 69068
rect 58676 69028 58682 69040
rect 60642 69028 60648 69040
rect 60700 69028 60706 69080
rect 69658 69028 69664 69080
rect 69716 69068 69722 69080
rect 71774 69068 71780 69080
rect 69716 69040 71780 69068
rect 69716 69028 69722 69040
rect 71774 69028 71780 69040
rect 71832 69028 71838 69080
rect 73062 69028 73068 69080
rect 73120 69068 73126 69080
rect 73890 69068 73896 69080
rect 73120 69040 73896 69068
rect 73120 69028 73126 69040
rect 73890 69028 73896 69040
rect 73948 69028 73954 69080
rect 75362 69028 75368 69080
rect 75420 69068 75426 69080
rect 75822 69068 75828 69080
rect 75420 69040 75828 69068
rect 75420 69028 75426 69040
rect 75822 69028 75828 69040
rect 75880 69028 75886 69080
rect 76742 69028 76748 69080
rect 76800 69068 76806 69080
rect 77202 69068 77208 69080
rect 76800 69040 77208 69068
rect 76800 69028 76806 69040
rect 77202 69028 77208 69040
rect 77260 69028 77266 69080
rect 77386 69028 77392 69080
rect 77444 69068 77450 69080
rect 79318 69068 79324 69080
rect 77444 69040 79324 69068
rect 77444 69028 77450 69040
rect 79318 69028 79324 69040
rect 79376 69028 79382 69080
rect 80238 69028 80244 69080
rect 80296 69068 80302 69080
rect 81342 69068 81348 69080
rect 80296 69040 81348 69068
rect 80296 69028 80302 69040
rect 81342 69028 81348 69040
rect 81400 69028 81406 69080
rect 82998 69028 83004 69080
rect 83056 69068 83062 69080
rect 84102 69068 84108 69080
rect 83056 69040 84108 69068
rect 83056 69028 83062 69040
rect 84102 69028 84108 69040
rect 84160 69028 84166 69080
rect 87598 69028 87604 69080
rect 87656 69068 87662 69080
rect 91370 69068 91376 69080
rect 87656 69040 91376 69068
rect 87656 69028 87662 69040
rect 91370 69028 91376 69040
rect 91428 69028 91434 69080
rect 94590 69028 94596 69080
rect 94648 69068 94654 69080
rect 96246 69068 96252 69080
rect 94648 69040 96252 69068
rect 94648 69028 94654 69040
rect 96246 69028 96252 69040
rect 96304 69028 96310 69080
rect 98638 69028 98644 69080
rect 98696 69068 98702 69080
rect 99742 69068 99748 69080
rect 98696 69040 99748 69068
rect 98696 69028 98702 69040
rect 99742 69028 99748 69040
rect 99800 69028 99806 69080
rect 103974 69028 103980 69080
rect 104032 69068 104038 69080
rect 104802 69068 104808 69080
rect 104032 69040 104808 69068
rect 104032 69028 104038 69040
rect 104802 69028 104808 69040
rect 104860 69028 104866 69080
rect 105354 69028 105360 69080
rect 105412 69068 105418 69080
rect 106090 69068 106096 69080
rect 105412 69040 106096 69068
rect 105412 69028 105418 69040
rect 106090 69028 106096 69040
rect 106148 69028 106154 69080
rect 125502 69028 125508 69080
rect 125560 69068 125566 69080
rect 128998 69068 129004 69080
rect 125560 69040 129004 69068
rect 125560 69028 125566 69040
rect 128998 69028 129004 69040
rect 129056 69028 129062 69080
rect 133782 69028 133788 69080
rect 133840 69068 133846 69080
rect 135346 69068 135352 69080
rect 133840 69040 135352 69068
rect 133840 69028 133846 69040
rect 135346 69028 135352 69040
rect 135404 69028 135410 69080
rect 136726 69028 136732 69080
rect 136784 69068 136790 69080
rect 137830 69068 137836 69080
rect 136784 69040 137836 69068
rect 136784 69028 136790 69040
rect 137830 69028 137836 69040
rect 137888 69028 137894 69080
rect 138106 69028 138112 69080
rect 138164 69068 138170 69080
rect 139302 69068 139308 69080
rect 138164 69040 139308 69068
rect 138164 69028 138170 69040
rect 139302 69028 139308 69040
rect 139360 69028 139366 69080
rect 139578 69028 139584 69080
rect 139636 69068 139642 69080
rect 140682 69068 140688 69080
rect 139636 69040 140688 69068
rect 139636 69028 139642 69040
rect 140682 69028 140688 69040
rect 140740 69028 140746 69080
rect 140958 69028 140964 69080
rect 141016 69068 141022 69080
rect 142062 69068 142068 69080
rect 141016 69040 142068 69068
rect 141016 69028 141022 69040
rect 142062 69028 142068 69040
rect 142120 69028 142126 69080
rect 142338 69028 142344 69080
rect 142396 69068 142402 69080
rect 143442 69068 143448 69080
rect 142396 69040 143448 69068
rect 142396 69028 142402 69040
rect 143442 69028 143448 69040
rect 143500 69028 143506 69080
rect 143718 69028 143724 69080
rect 143776 69068 143782 69080
rect 144638 69068 144644 69080
rect 143776 69040 144644 69068
rect 143776 69028 143782 69040
rect 144638 69028 144644 69040
rect 144696 69028 144702 69080
rect 145098 69028 145104 69080
rect 145156 69068 145162 69080
rect 146110 69068 146116 69080
rect 145156 69040 146116 69068
rect 145156 69028 145162 69040
rect 146110 69028 146116 69040
rect 146168 69028 146174 69080
rect 146478 69028 146484 69080
rect 146536 69068 146542 69080
rect 147582 69068 147588 69080
rect 146536 69040 147588 69068
rect 146536 69028 146542 69040
rect 147582 69028 147588 69040
rect 147640 69028 147646 69080
rect 147950 69028 147956 69080
rect 148008 69068 148014 69080
rect 148870 69068 148876 69080
rect 148008 69040 148876 69068
rect 148008 69028 148014 69040
rect 148870 69028 148876 69040
rect 148928 69028 148934 69080
rect 149330 69028 149336 69080
rect 149388 69068 149394 69080
rect 150250 69068 150256 69080
rect 149388 69040 150256 69068
rect 149388 69028 149394 69040
rect 150250 69028 150256 69040
rect 150308 69028 150314 69080
rect 150710 69028 150716 69080
rect 150768 69068 150774 69080
rect 151722 69068 151728 69080
rect 150768 69040 151728 69068
rect 150768 69028 150774 69040
rect 151722 69028 151728 69040
rect 151780 69028 151786 69080
rect 152090 69028 152096 69080
rect 152148 69068 152154 69080
rect 153010 69068 153016 69080
rect 152148 69040 153016 69068
rect 152148 69028 152154 69040
rect 153010 69028 153016 69040
rect 153068 69028 153074 69080
rect 153470 69028 153476 69080
rect 153528 69068 153534 69080
rect 154482 69068 154488 69080
rect 153528 69040 154488 69068
rect 153528 69028 153534 69040
rect 154482 69028 154488 69040
rect 154540 69028 154546 69080
rect 159082 69028 159088 69080
rect 159140 69068 159146 69080
rect 159910 69068 159916 69080
rect 159140 69040 159916 69068
rect 159140 69028 159146 69040
rect 159910 69028 159916 69040
rect 159968 69028 159974 69080
rect 160462 69028 160468 69080
rect 160520 69068 160526 69080
rect 161382 69068 161388 69080
rect 160520 69040 161388 69068
rect 160520 69028 160526 69040
rect 161382 69028 161388 69040
rect 161440 69028 161446 69080
rect 161842 69028 161848 69080
rect 161900 69068 161906 69080
rect 162670 69068 162676 69080
rect 161900 69040 162676 69068
rect 161900 69028 161906 69040
rect 162670 69028 162676 69040
rect 162728 69028 162734 69080
rect 166074 69028 166080 69080
rect 166132 69068 166138 69080
rect 166810 69068 166816 69080
rect 166132 69040 166816 69068
rect 166132 69028 166138 69040
rect 166810 69028 166816 69040
rect 166868 69028 166874 69080
rect 167454 69028 167460 69080
rect 167512 69068 167518 69080
rect 168282 69068 168288 69080
rect 167512 69040 168288 69068
rect 167512 69028 167518 69040
rect 168282 69028 168288 69040
rect 168340 69028 168346 69080
rect 168834 69028 168840 69080
rect 168892 69068 168898 69080
rect 169662 69068 169668 69080
rect 168892 69040 169668 69068
rect 168892 69028 168898 69040
rect 169662 69028 169668 69040
rect 169720 69028 169726 69080
rect 170214 69028 170220 69080
rect 170272 69068 170278 69080
rect 170950 69068 170956 69080
rect 170272 69040 170956 69068
rect 170272 69028 170278 69040
rect 170950 69028 170956 69040
rect 171008 69028 171014 69080
rect 171594 69028 171600 69080
rect 171652 69068 171658 69080
rect 173158 69068 173164 69080
rect 171652 69040 173164 69068
rect 171652 69028 171658 69040
rect 173158 69028 173164 69040
rect 173216 69028 173222 69080
rect 174446 69028 174452 69080
rect 174504 69068 174510 69080
rect 175090 69068 175096 69080
rect 174504 69040 175096 69068
rect 174504 69028 174510 69040
rect 175090 69028 175096 69040
rect 175148 69028 175154 69080
rect 175826 69028 175832 69080
rect 175884 69068 175890 69080
rect 176470 69068 176476 69080
rect 175884 69040 176476 69068
rect 175884 69028 175890 69040
rect 176470 69028 176476 69040
rect 176528 69028 176534 69080
rect 178586 69028 178592 69080
rect 178644 69068 178650 69080
rect 179230 69068 179236 69080
rect 178644 69040 179236 69068
rect 178644 69028 178650 69040
rect 179230 69028 179236 69040
rect 179288 69028 179294 69080
rect 179966 69028 179972 69080
rect 180024 69068 180030 69080
rect 180610 69068 180616 69080
rect 180024 69040 180616 69068
rect 180024 69028 180030 69040
rect 180610 69028 180616 69040
rect 180668 69028 180674 69080
rect 181438 69028 181444 69080
rect 181496 69068 181502 69080
rect 182082 69068 182088 69080
rect 181496 69040 182088 69068
rect 181496 69028 181502 69040
rect 182082 69028 182088 69040
rect 182140 69028 182146 69080
rect 182818 69028 182824 69080
rect 182876 69068 182882 69080
rect 183370 69068 183376 69080
rect 182876 69040 183376 69068
rect 182876 69028 182882 69040
rect 183370 69028 183376 69040
rect 183428 69028 183434 69080
rect 184198 69028 184204 69080
rect 184256 69068 184262 69080
rect 184842 69068 184848 69080
rect 184256 69040 184848 69068
rect 184256 69028 184262 69040
rect 184842 69028 184848 69040
rect 184900 69028 184906 69080
rect 185578 69028 185584 69080
rect 185636 69068 185642 69080
rect 186222 69068 186228 69080
rect 185636 69040 186228 69068
rect 185636 69028 185642 69040
rect 186222 69028 186228 69040
rect 186280 69028 186286 69080
rect 186958 69028 186964 69080
rect 187016 69068 187022 69080
rect 187510 69068 187516 69080
rect 187016 69040 187516 69068
rect 187016 69028 187022 69040
rect 187510 69028 187516 69040
rect 187568 69028 187574 69080
rect 188338 69028 188344 69080
rect 188396 69068 188402 69080
rect 188982 69068 188988 69080
rect 188396 69040 188988 69068
rect 188396 69028 188402 69040
rect 188982 69028 188988 69040
rect 189040 69028 189046 69080
rect 189810 69028 189816 69080
rect 189868 69068 189874 69080
rect 190362 69068 190368 69080
rect 189868 69040 190368 69068
rect 189868 69028 189874 69040
rect 190362 69028 190368 69040
rect 190420 69028 190426 69080
rect 191190 69028 191196 69080
rect 191248 69068 191254 69080
rect 191742 69068 191748 69080
rect 191248 69040 191748 69068
rect 191248 69028 191254 69040
rect 191742 69028 191748 69040
rect 191800 69028 191806 69080
rect 191834 69028 191840 69080
rect 191892 69068 191898 69080
rect 193122 69068 193128 69080
rect 191892 69040 193128 69068
rect 191892 69028 191898 69040
rect 193122 69028 193128 69040
rect 193180 69028 193186 69080
rect 195330 69028 195336 69080
rect 195388 69068 195394 69080
rect 195790 69068 195796 69080
rect 195388 69040 195796 69068
rect 195388 69028 195394 69040
rect 195790 69028 195796 69040
rect 195848 69028 195854 69080
rect 196710 69028 196716 69080
rect 196768 69068 196774 69080
rect 197262 69068 197268 69080
rect 196768 69040 197268 69068
rect 196768 69028 196774 69040
rect 197262 69028 197268 69040
rect 197320 69028 197326 69080
rect 198182 69028 198188 69080
rect 198240 69068 198246 69080
rect 198642 69068 198648 69080
rect 198240 69040 198648 69068
rect 198240 69028 198246 69040
rect 198642 69028 198648 69040
rect 198700 69028 198706 69080
rect 199562 69028 199568 69080
rect 199620 69068 199626 69080
rect 200022 69068 200028 69080
rect 199620 69040 200028 69068
rect 199620 69028 199626 69040
rect 200022 69028 200028 69040
rect 200080 69028 200086 69080
rect 200206 69028 200212 69080
rect 200264 69068 200270 69080
rect 201402 69068 201408 69080
rect 200264 69040 201408 69068
rect 200264 69028 200270 69040
rect 201402 69028 201408 69040
rect 201460 69028 201466 69080
rect 201678 69028 201684 69080
rect 201736 69068 201742 69080
rect 202782 69068 202788 69080
rect 201736 69040 202788 69068
rect 201736 69028 201742 69040
rect 202782 69028 202788 69040
rect 202840 69028 202846 69080
rect 203058 69028 203064 69080
rect 203116 69068 203122 69080
rect 204162 69068 204168 69080
rect 203116 69040 204168 69068
rect 203116 69028 203122 69040
rect 204162 69028 204168 69040
rect 204220 69028 204226 69080
rect 206756 69068 206784 69108
rect 207934 69096 207940 69148
rect 207992 69136 207998 69148
<<<<<<< HEAD
rect 213546 69136 213552 69148
rect 207992 69108 213552 69136
rect 207992 69096 207998 69108
rect 213546 69096 213552 69108
rect 213604 69096 213610 69148
=======
rect 213638 69136 213644 69148
rect 207992 69108 213644 69136
rect 207992 69096 207998 69108
rect 213638 69096 213644 69108
rect 213696 69096 213702 69148
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 248414 69096 248420 69148
rect 248472 69136 248478 69148
rect 249702 69136 249708 69148
rect 248472 69108 249708 69136
rect 248472 69096 248478 69108
rect 249702 69096 249708 69108
rect 249760 69096 249766 69148
rect 251174 69096 251180 69148
rect 251232 69136 251238 69148
rect 252462 69136 252468 69148
rect 251232 69108 252468 69136
rect 251232 69096 251238 69108
rect 252462 69096 252468 69108
rect 252520 69096 252526 69148
rect 252554 69096 252560 69148
rect 252612 69136 252618 69148
rect 253842 69136 253848 69148
rect 252612 69108 253848 69136
rect 252612 69096 252618 69108
rect 253842 69096 253848 69108
rect 253900 69096 253906 69148
rect 253934 69096 253940 69148
rect 253992 69136 253998 69148
rect 255222 69136 255228 69148
rect 253992 69108 255228 69136
rect 253992 69096 253998 69108
rect 255222 69096 255228 69108
rect 255280 69096 255286 69148
rect 255406 69096 255412 69148
rect 255464 69136 255470 69148
rect 256602 69136 256608 69148
rect 255464 69108 256608 69136
rect 255464 69096 255470 69108
rect 256602 69096 256608 69108
rect 256660 69096 256666 69148
rect 256786 69096 256792 69148
rect 256844 69136 256850 69148
rect 257890 69136 257896 69148
rect 256844 69108 257896 69136
rect 256844 69096 256850 69108
rect 257890 69096 257896 69108
rect 257948 69096 257954 69148
rect 258166 69096 258172 69148
rect 258224 69136 258230 69148
rect 259270 69136 259276 69148
rect 258224 69108 259276 69136
rect 258224 69096 258230 69108
rect 259270 69096 259276 69108
rect 259328 69096 259334 69148
rect 260926 69096 260932 69148
rect 260984 69136 260990 69148
rect 262030 69136 262036 69148
rect 260984 69108 262036 69136
rect 260984 69096 260990 69108
rect 262030 69096 262036 69108
rect 262088 69096 262094 69148
rect 262306 69096 262312 69148
rect 262364 69136 262370 69148
rect 263410 69136 263416 69148
rect 262364 69108 263416 69136
rect 262364 69096 262370 69108
rect 263410 69096 263416 69108
rect 263468 69096 263474 69148
rect 310514 69096 310520 69148
rect 310572 69136 310578 69148
rect 311802 69136 311808 69148
rect 310572 69108 311808 69136
rect 310572 69096 310578 69108
rect 311802 69096 311808 69108
rect 311860 69096 311866 69148
rect 327718 69096 327724 69148
rect 327776 69136 327782 69148
rect 332778 69136 332784 69148
rect 327776 69108 332784 69136
rect 327776 69096 327782 69108
rect 332778 69096 332784 69108
rect 332836 69096 332842 69148
rect 389358 69096 389364 69148
rect 389416 69136 389422 69148
rect 390370 69136 390376 69148
rect 389416 69108 390376 69136
rect 389416 69096 389422 69108
rect 390370 69096 390376 69108
rect 390428 69096 390434 69148
<<<<<<< HEAD
rect 390738 69096 390744 69148
rect 390796 69136 390802 69148
rect 392394 69136 392400 69148
rect 390796 69108 392400 69136
rect 390796 69096 390802 69108
rect 392394 69096 392400 69108
rect 392452 69096 392458 69148
rect 403342 69096 403348 69148
rect 403400 69136 403406 69148
rect 404170 69136 404176 69148
rect 403400 69108 404176 69136
rect 403400 69096 403406 69108
rect 404170 69096 404176 69108
rect 404228 69096 404234 69148
=======
rect 401870 69096 401876 69148
rect 401928 69136 401934 69148
rect 403710 69136 403716 69148
rect 401928 69108 403716 69136
rect 401928 69096 401934 69108
rect 403710 69096 403716 69108
rect 403768 69096 403774 69148
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 209961 69071 210019 69077
rect 209961 69068 209973 69071
rect 206756 69040 209973 69068
rect 209961 69037 209973 69040
rect 210007 69037 210019 69071
rect 209961 69031 210019 69037
rect 210050 69028 210056 69080
rect 210108 69068 210114 69080
rect 210970 69068 210976 69080
rect 210108 69040 210976 69068
rect 210108 69028 210114 69040
rect 210970 69028 210976 69040
rect 211028 69028 211034 69080
rect 211430 69028 211436 69080
rect 211488 69068 211494 69080
rect 212350 69068 212356 69080
rect 211488 69040 212356 69068
rect 211488 69028 211494 69040
rect 212350 69028 212356 69040
rect 212408 69028 212414 69080
rect 212810 69028 212816 69080
rect 212868 69068 212874 69080
rect 213822 69068 213828 69080
rect 212868 69040 213828 69068
rect 212868 69028 212874 69040
rect 213822 69028 213828 69040
rect 213880 69028 213886 69080
rect 214190 69028 214196 69080
rect 214248 69068 214254 69080
rect 215110 69068 215116 69080
rect 214248 69040 215116 69068
rect 214248 69028 214254 69040
rect 215110 69028 215116 69040
rect 215168 69028 215174 69080
rect 215570 69028 215576 69080
rect 215628 69068 215634 69080
rect 216490 69068 216496 69080
rect 215628 69040 216496 69068
rect 215628 69028 215634 69040
rect 216490 69028 216496 69040
rect 216548 69028 216554 69080
rect 216950 69028 216956 69080
rect 217008 69068 217014 69080
rect 217870 69068 217876 69080
rect 217008 69040 217876 69068
rect 217008 69028 217014 69040
rect 217870 69028 217876 69040
rect 217928 69028 217934 69080
rect 218422 69028 218428 69080
rect 218480 69068 218486 69080
rect 218974 69068 218980 69080
rect 218480 69040 218980 69068
rect 218480 69028 218486 69040
rect 218974 69028 218980 69040
rect 219032 69028 219038 69080
rect 219802 69028 219808 69080
rect 219860 69068 219866 69080
rect 220630 69068 220636 69080
rect 219860 69040 220636 69068
rect 219860 69028 219866 69040
rect 220630 69028 220636 69040
rect 220688 69028 220694 69080
rect 221182 69028 221188 69080
rect 221240 69068 221246 69080
rect 222102 69068 222108 69080
rect 221240 69040 222108 69068
rect 221240 69028 221246 69040
rect 222102 69028 222108 69040
rect 222160 69028 222166 69080
rect 232498 69028 232504 69080
rect 232556 69068 232562 69080
rect 235074 69068 235080 69080
rect 232556 69040 235080 69068
rect 232556 69028 232562 69040
rect 235074 69028 235080 69040
rect 235132 69028 235138 69080
rect 242158 69028 242164 69080
rect 242216 69068 242222 69080
rect 243446 69068 243452 69080
rect 242216 69040 243452 69068
rect 242216 69028 242222 69040
rect 243446 69028 243452 69040
rect 243504 69028 243510 69080
rect 249058 69028 249064 69080
rect 249116 69068 249122 69080
rect 249610 69068 249616 69080
rect 249116 69040 249616 69068
rect 249116 69028 249122 69040
rect 249610 69028 249616 69040
rect 249668 69028 249674 69080
rect 249794 69028 249800 69080
rect 249852 69068 249858 69080
rect 251082 69068 251088 69080
rect 249852 69040 251088 69068
rect 249852 69028 249858 69040
rect 251082 69028 251088 69040
rect 251140 69028 251146 69080
rect 251910 69028 251916 69080
rect 251968 69068 251974 69080
rect 252370 69068 252376 69080
rect 251968 69040 252376 69068
rect 251968 69028 251974 69040
rect 252370 69028 252376 69040
rect 252428 69028 252434 69080
rect 253290 69028 253296 69080
rect 253348 69068 253354 69080
rect 253750 69068 253756 69080
rect 253348 69040 253756 69068
rect 253348 69028 253354 69040
rect 253750 69028 253756 69040
rect 253808 69028 253814 69080
rect 254670 69028 254676 69080
rect 254728 69068 254734 69080
rect 255130 69068 255136 69080
rect 254728 69040 255136 69068
rect 254728 69028 254734 69040
rect 255130 69028 255136 69040
rect 255188 69028 255194 69080
rect 256050 69028 256056 69080
rect 256108 69068 256114 69080
rect 256510 69068 256516 69080
rect 256108 69040 256516 69068
rect 256108 69028 256114 69040
rect 256510 69028 256516 69040
rect 256568 69028 256574 69080
rect 257430 69028 257436 69080
rect 257488 69068 257494 69080
rect 257982 69068 257988 69080
rect 257488 69040 257988 69068
rect 257488 69028 257494 69040
rect 257982 69028 257988 69040
rect 258040 69028 258046 69080
rect 258902 69028 258908 69080
rect 258960 69068 258966 69080
rect 259362 69068 259368 69080
rect 258960 69040 259368 69068
rect 258960 69028 258966 69040
rect 259362 69028 259368 69040
rect 259420 69028 259426 69080
rect 259546 69028 259552 69080
rect 259604 69068 259610 69080
rect 260742 69068 260748 69080
rect 259604 69040 260748 69068
rect 259604 69028 259610 69040
rect 260742 69028 260748 69040
rect 260800 69028 260806 69080
rect 261662 69028 261668 69080
rect 261720 69068 261726 69080
rect 262122 69068 262128 69080
rect 261720 69040 262128 69068
rect 261720 69028 261726 69040
rect 262122 69028 262128 69040
rect 262180 69028 262186 69080
rect 263042 69028 263048 69080
rect 263100 69068 263106 69080
rect 263502 69068 263508 69080
rect 263100 69040 263508 69068
rect 263100 69028 263106 69040
rect 263502 69028 263508 69040
rect 263560 69028 263566 69080
rect 263778 69028 263784 69080
rect 263836 69068 263842 69080
rect 264882 69068 264888 69080
rect 263836 69040 264888 69068
rect 263836 69028 263842 69040
rect 264882 69028 264888 69040
rect 264940 69028 264946 69080
rect 265158 69028 265164 69080
rect 265216 69068 265222 69080
rect 266262 69068 266268 69080
rect 265216 69040 266268 69068
rect 265216 69028 265222 69040
rect 266262 69028 266268 69040
rect 266320 69028 266326 69080
rect 266538 69028 266544 69080
rect 266596 69068 266602 69080
rect 267642 69068 267648 69080
rect 266596 69040 267648 69068
rect 266596 69028 266602 69040
rect 267642 69028 267648 69040
rect 267700 69028 267706 69080
rect 267918 69028 267924 69080
rect 267976 69068 267982 69080
rect 269022 69068 269028 69080
rect 267976 69040 269028 69068
rect 267976 69028 267982 69040
rect 269022 69028 269028 69040
rect 269080 69028 269086 69080
rect 269298 69028 269304 69080
rect 269356 69068 269362 69080
rect 270310 69068 270316 69080
rect 269356 69040 270316 69068
rect 269356 69028 269362 69040
rect 270310 69028 270316 69040
rect 270368 69028 270374 69080
rect 270678 69028 270684 69080
rect 270736 69068 270742 69080
rect 271690 69068 271696 69080
rect 270736 69040 271696 69068
rect 270736 69028 270742 69040
rect 271690 69028 271696 69040
rect 271748 69028 271754 69080
rect 273530 69028 273536 69080
rect 273588 69068 273594 69080
rect 274450 69068 274456 69080
rect 273588 69040 274456 69068
rect 273588 69028 273594 69040
rect 274450 69028 274456 69040
rect 274508 69028 274514 69080
rect 274910 69028 274916 69080
rect 274968 69068 274974 69080
rect 275830 69068 275836 69080
rect 274968 69040 275836 69068
rect 274968 69028 274974 69040
rect 275830 69028 275836 69040
rect 275888 69028 275894 69080
rect 276290 69028 276296 69080
rect 276348 69068 276354 69080
rect 277210 69068 277216 69080
rect 276348 69040 277216 69068
rect 276348 69028 276354 69040
rect 277210 69028 277216 69040
rect 277268 69028 277274 69080
rect 277670 69028 277676 69080
rect 277728 69068 277734 69080
rect 278590 69068 278596 69080
rect 277728 69040 278596 69068
rect 277728 69028 277734 69040
rect 278590 69028 278596 69040
rect 278648 69028 278654 69080
rect 279050 69028 279056 69080
rect 279108 69068 279114 69080
rect 279970 69068 279976 69080
rect 279108 69040 279976 69068
rect 279108 69028 279114 69040
rect 279970 69028 279976 69040
rect 280028 69028 280034 69080
rect 280522 69028 280528 69080
rect 280580 69068 280586 69080
rect 281350 69068 281356 69080
rect 280580 69040 281356 69068
rect 280580 69028 280586 69040
rect 281350 69028 281356 69040
rect 281408 69028 281414 69080
rect 281902 69028 281908 69080
rect 281960 69068 281966 69080
rect 282730 69068 282736 69080
rect 281960 69040 282736 69068
rect 281960 69028 281966 69040
rect 282730 69028 282736 69040
rect 282788 69028 282794 69080
rect 283282 69028 283288 69080
rect 283340 69068 283346 69080
rect 284202 69068 284208 69080
rect 283340 69040 284208 69068
rect 283340 69028 283346 69040
rect 284202 69028 284208 69040
rect 284260 69028 284266 69080
rect 284662 69028 284668 69080
rect 284720 69068 284726 69080
rect 285490 69068 285496 69080
rect 284720 69040 285496 69068
rect 284720 69028 284726 69040
rect 285490 69028 285496 69040
rect 285548 69028 285554 69080
rect 286042 69028 286048 69080
rect 286100 69068 286106 69080
rect 286870 69068 286876 69080
rect 286100 69040 286876 69068
rect 286100 69028 286106 69040
rect 286870 69028 286876 69040
rect 286928 69028 286934 69080
rect 287422 69028 287428 69080
rect 287480 69068 287486 69080
rect 288342 69068 288348 69080
rect 287480 69040 288348 69068
rect 287480 69028 287486 69040
rect 288342 69028 288348 69040
rect 288400 69028 288406 69080
rect 288894 69028 288900 69080
rect 288952 69068 288958 69080
rect 289722 69068 289728 69080
rect 288952 69040 289728 69068
rect 288952 69028 288958 69040
rect 289722 69028 289728 69040
rect 289780 69028 289786 69080
rect 290918 69028 290924 69080
rect 290976 69068 290982 69080
rect 293770 69068 293776 69080
rect 290976 69040 293776 69068
rect 290976 69028 290982 69040
rect 293770 69028 293776 69040
rect 293828 69028 293834 69080
rect 297266 69028 297272 69080
rect 297324 69068 297330 69080
rect 298002 69068 298008 69080
rect 297324 69040 298008 69068
rect 297324 69028 297330 69040
rect 298002 69028 298008 69040
rect 298060 69028 298066 69080
rect 298646 69028 298652 69080
rect 298704 69068 298710 69080
rect 299290 69068 299296 69080
rect 298704 69040 299296 69068
rect 298704 69028 298710 69040
rect 299290 69028 299296 69040
rect 299348 69028 299354 69080
rect 300026 69028 300032 69080
rect 300084 69068 300090 69080
rect 300670 69068 300676 69080
rect 300084 69040 300676 69068
rect 300084 69028 300090 69040
rect 300670 69028 300676 69040
rect 300728 69028 300734 69080
rect 301406 69028 301412 69080
rect 301464 69068 301470 69080
rect 302142 69068 302148 69080
rect 301464 69040 302148 69068
rect 301464 69028 301470 69040
rect 302142 69028 302148 69040
rect 302200 69028 302206 69080
rect 302786 69028 302792 69080
rect 302844 69068 302850 69080
rect 303522 69068 303528 69080
rect 302844 69040 303528 69068
rect 302844 69028 302850 69040
rect 303522 69028 303528 69040
rect 303580 69028 303586 69080
rect 304258 69028 304264 69080
rect 304316 69068 304322 69080
rect 304810 69068 304816 69080
rect 304316 69040 304816 69068
rect 304316 69028 304322 69040
rect 304810 69028 304816 69040
rect 304868 69028 304874 69080
rect 305638 69028 305644 69080
rect 305696 69068 305702 69080
rect 306190 69068 306196 69080
rect 305696 69040 306196 69068
rect 305696 69028 305702 69040
rect 306190 69028 306196 69040
rect 306248 69028 306254 69080
rect 307018 69028 307024 69080
rect 307076 69068 307082 69080
rect 307662 69068 307668 69080
rect 307076 69040 307668 69068
rect 307076 69028 307082 69040
rect 307662 69028 307668 69040
rect 307720 69028 307726 69080
rect 308398 69028 308404 69080
rect 308456 69068 308462 69080
rect 309042 69068 309048 69080
rect 308456 69040 309048 69068
rect 308456 69028 308462 69040
rect 309042 69028 309048 69040
rect 309100 69028 309106 69080
rect 309778 69028 309784 69080
rect 309836 69068 309842 69080
rect 310422 69068 310428 69080
rect 309836 69040 310428 69068
rect 309836 69028 309842 69040
rect 310422 69028 310428 69040
rect 310480 69028 310486 69080
rect 311158 69028 311164 69080
rect 311216 69068 311222 69080
rect 311710 69068 311716 69080
rect 311216 69040 311716 69068
rect 311216 69028 311222 69040
rect 311710 69028 311716 69040
rect 311768 69028 311774 69080
rect 311894 69028 311900 69080
rect 311952 69068 311958 69080
rect 313090 69068 313096 69080
rect 311952 69040 313096 69068
rect 311952 69028 311958 69040
rect 313090 69028 313096 69040
rect 313148 69028 313154 69080
rect 331858 69028 331864 69080
rect 331916 69068 331922 69080
rect 333514 69068 333520 69080
rect 331916 69040 333520 69068
rect 331916 69028 331922 69040
rect 333514 69028 333520 69040
rect 333572 69028 333578 69080
rect 359366 69028 359372 69080
rect 359424 69068 359430 69080
rect 360102 69068 360108 69080
rect 359424 69040 360108 69068
rect 359424 69028 359430 69040
rect 360102 69028 360108 69040
rect 360160 69028 360166 69080
rect 360746 69028 360752 69080
rect 360804 69068 360810 69080
rect 361390 69068 361396 69080
rect 360804 69040 361396 69068
rect 360804 69028 360810 69040
rect 361390 69028 361396 69040
rect 361448 69028 361454 69080
rect 362126 69028 362132 69080
rect 362184 69068 362190 69080
rect 362862 69068 362868 69080
rect 362184 69040 362868 69068
rect 362184 69028 362190 69040
rect 362862 69028 362868 69040
rect 362920 69028 362926 69080
rect 363506 69028 363512 69080
rect 363564 69068 363570 69080
rect 364242 69068 364248 69080
rect 363564 69040 364248 69068
rect 363564 69028 363570 69040
rect 364242 69028 364248 69040
rect 364300 69028 364306 69080
rect 364886 69028 364892 69080
rect 364944 69068 364950 69080
rect 365622 69068 365628 69080
rect 364944 69040 365628 69068
rect 364944 69028 364950 69040
rect 365622 69028 365628 69040
rect 365680 69028 365686 69080
rect 366358 69028 366364 69080
rect 366416 69068 366422 69080
rect 366910 69068 366916 69080
rect 366416 69040 366916 69068
rect 366416 69028 366422 69040
rect 366910 69028 366916 69040
rect 366968 69028 366974 69080
rect 369118 69028 369124 69080
rect 369176 69068 369182 69080
rect 369670 69068 369676 69080
rect 369176 69040 369676 69068
rect 369176 69028 369182 69040
rect 369670 69028 369676 69040
rect 369728 69028 369734 69080
rect 373258 69028 373264 69080
rect 373316 69068 373322 69080
rect 373902 69068 373908 69080
rect 373316 69040 373908 69068
rect 373316 69028 373322 69040
rect 373902 69028 373908 69040
rect 373960 69028 373966 69080
rect 374730 69028 374736 69080
rect 374788 69068 374794 69080
rect 375282 69068 375288 69080
rect 374788 69040 375288 69068
rect 374788 69028 374794 69040
rect 375282 69028 375288 69040
rect 375340 69028 375346 69080
rect 376110 69028 376116 69080
rect 376168 69068 376174 69080
rect 376662 69068 376668 69080
rect 376168 69040 376668 69068
rect 376168 69028 376174 69040
rect 376662 69028 376668 69040
rect 376720 69028 376726 69080
rect 377490 69028 377496 69080
rect 377548 69068 377554 69080
rect 378042 69068 378048 69080
rect 377548 69040 378048 69068
rect 377548 69028 377554 69040
rect 378042 69028 378048 69040
rect 378100 69028 378106 69080
rect 378870 69028 378876 69080
rect 378928 69068 378934 69080
rect 379422 69068 379428 69080
rect 378928 69040 379428 69068
rect 378928 69028 378934 69040
rect 379422 69028 379428 69040
rect 379480 69028 379486 69080
rect 380250 69028 380256 69080
rect 380308 69068 380314 69080
rect 380802 69068 380808 69080
rect 380308 69040 380808 69068
rect 380308 69028 380314 69040
rect 380802 69028 380808 69040
rect 380860 69028 380866 69080
rect 381630 69028 381636 69080
rect 381688 69068 381694 69080
rect 382182 69068 382188 69080
rect 381688 69040 382188 69068
rect 381688 69028 381694 69040
rect 382182 69028 382188 69040
rect 382240 69028 382246 69080
rect 382366 69028 382372 69080
rect 382424 69068 382430 69080
rect 383562 69068 383568 69080
rect 382424 69040 383568 69068
rect 382424 69028 382430 69040
rect 383562 69028 383568 69040
rect 383620 69028 383626 69080
rect 385862 69028 385868 69080
rect 385920 69068 385926 69080
rect 386322 69068 386328 69080
rect 385920 69040 386328 69068
rect 385920 69028 385926 69040
rect 386322 69028 386328 69040
rect 386380 69028 386386 69080
rect 388622 69028 388628 69080
rect 388680 69068 388686 69080
rect 389082 69068 389088 69080
rect 388680 69040 389088 69068
rect 388680 69028 388686 69040
rect 389082 69028 389088 69040
rect 389140 69028 389146 69080
rect 390002 69028 390008 69080
rect 390060 69068 390066 69080
rect 390462 69068 390468 69080
rect 390060 69040 390468 69068
rect 390060 69028 390066 69040
rect 390462 69028 390468 69040
rect 390520 69028 390526 69080
<<<<<<< HEAD
=======
rect 390738 69028 390744 69080
rect 390796 69068 390802 69080
rect 391934 69068 391940 69080
rect 390796 69040 391940 69068
rect 390796 69028 390802 69040
rect 391934 69028 391940 69040
rect 391992 69028 391998 69080
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 392118 69028 392124 69080
rect 392176 69068 392182 69080
rect 393130 69068 393136 69080
rect 392176 69040 393136 69068
rect 392176 69028 392182 69040
rect 393130 69028 393136 69040
rect 393188 69028 393194 69080
rect 393498 69028 393504 69080
rect 393556 69068 393562 69080
rect 394510 69068 394516 69080
rect 393556 69040 394516 69068
rect 393556 69028 393562 69040
rect 394510 69028 394516 69040
rect 394568 69028 394574 69080
rect 394970 69028 394976 69080
rect 395028 69068 395034 69080
rect 395890 69068 395896 69080
rect 395028 69040 395896 69068
rect 395028 69028 395034 69040
rect 395890 69028 395896 69040
rect 395948 69028 395954 69080
rect 396350 69028 396356 69080
rect 396408 69068 396414 69080
rect 397270 69068 397276 69080
rect 396408 69040 397276 69068
rect 396408 69028 396414 69040
rect 397270 69028 397276 69040
rect 397328 69028 397334 69080
rect 397730 69028 397736 69080
rect 397788 69068 397794 69080
rect 398742 69068 398748 69080
rect 397788 69040 398748 69068
rect 397788 69028 397794 69040
rect 398742 69028 398748 69040
rect 398800 69028 398806 69080
rect 399110 69028 399116 69080
rect 399168 69068 399174 69080
rect 400122 69068 400128 69080
rect 399168 69040 400128 69068
rect 399168 69028 399174 69040
rect 400122 69028 400128 69040
rect 400180 69028 400186 69080
rect 400490 69028 400496 69080
rect 400548 69068 400554 69080
rect 401502 69068 401508 69080
rect 400548 69040 401508 69068
rect 400548 69028 400554 69040
rect 401502 69028 401508 69040
rect 401560 69028 401566 69080
<<<<<<< HEAD
rect 401870 69028 401876 69080
rect 401928 69068 401934 69080
rect 404262 69068 404268 69080
rect 401928 69040 404268 69068
rect 401928 69028 401934 69040
=======
rect 403342 69028 403348 69080
rect 403400 69068 403406 69080
rect 404262 69068 404268 69080
rect 403400 69040 404268 69068
rect 403400 69028 403406 69040
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 404262 69028 404268 69040
rect 404320 69028 404326 69080
rect 384482 68824 384488 68876
rect 384540 68864 384546 68876
rect 492674 68864 492680 68876
rect 384540 68836 492680 68864
rect 384540 68824 384546 68836
rect 492674 68824 492680 68836
rect 492732 68824 492738 68876
rect 55122 68756 55128 68808
rect 55180 68796 55186 68808
rect 70394 68796 70400 68808
rect 55180 68768 70400 68796
rect 55180 68756 55186 68768
rect 70394 68756 70400 68768
rect 70452 68756 70458 68808
rect 172330 68756 172336 68808
rect 172388 68796 172394 68808
rect 320174 68796 320180 68808
rect 172388 68768 320180 68796
rect 172388 68756 172394 68768
rect 320174 68756 320180 68768
rect 320232 68756 320238 68808
rect 386598 68756 386604 68808
rect 386656 68796 386662 68808
rect 503714 68796 503720 68808
rect 386656 68768 503720 68796
rect 386656 68756 386662 68768
rect 503714 68756 503720 68768
rect 503772 68756 503778 68808
rect 48222 68688 48228 68740
rect 48280 68728 48286 68740
rect 69014 68728 69020 68740
rect 48280 68700 69020 68728
rect 48280 68688 48286 68700
rect 69014 68688 69020 68700
rect 69072 68688 69078 68740
rect 177206 68688 177212 68740
rect 177264 68728 177270 68740
rect 345014 68728 345020 68740
rect 177264 68700 345020 68728
rect 177264 68688 177270 68700
rect 345014 68688 345020 68700
rect 345072 68688 345078 68740
rect 391474 68688 391480 68740
rect 391532 68728 391538 68740
rect 528554 68728 528560 68740
rect 391532 68700 528560 68728
rect 391532 68688 391538 68700
rect 528554 68688 528560 68700
rect 528612 68688 528618 68740
rect 37182 68620 37188 68672
rect 37240 68660 37246 68672
rect 65886 68660 65892 68672
rect 37240 68632 65892 68660
rect 37240 68620 37246 68632
rect 65886 68620 65892 68632
rect 65944 68620 65950 68672
rect 310330 68620 310336 68672
rect 310388 68660 310394 68672
rect 481634 68660 481640 68672
rect 310388 68632 481640 68660
rect 310388 68620 310394 68632
rect 481634 68620 481640 68632
rect 481692 68620 481698 68672
rect 14458 68552 14464 68604
rect 14516 68592 14522 68604
rect 62758 68592 62764 68604
rect 14516 68564 62764 68592
rect 14516 68552 14522 68564
rect 62758 68552 62764 68564
rect 62816 68552 62822 68604
<<<<<<< HEAD
rect 177298 68552 177304 68604
rect 177356 68592 177362 68604
rect 229554 68592 229560 68604
rect 177356 68564 229560 68592
rect 177356 68552 177362 68564
rect 229554 68552 229560 68564
rect 229612 68552 229618 68604
rect 244366 68552 244372 68604
rect 244424 68592 244430 68604
rect 245562 68592 245568 68604
rect 244424 68564 245568 68592
rect 244424 68552 244430 68564
rect 245562 68552 245568 68564
rect 245620 68552 245626 68604
rect 295886 68552 295892 68604
rect 295944 68592 295950 68604
rect 488534 68592 488540 68604
rect 295944 68564 488540 68592
rect 295944 68552 295950 68564
rect 488534 68552 488540 68564
rect 488592 68552 488598 68604
=======
rect 134518 68552 134524 68604
rect 134576 68592 134582 68604
rect 312538 68592 312544 68604
rect 134576 68564 312544 68592
rect 134576 68552 134582 68564
rect 312538 68552 312544 68564
rect 312596 68552 312602 68604
rect 314746 68552 314752 68604
rect 314804 68592 314810 68604
rect 315298 68592 315304 68604
rect 314804 68564 315304 68592
rect 314804 68552 314810 68564
rect 315298 68552 315304 68564
rect 315356 68552 315362 68604
rect 403710 68552 403716 68604
rect 403768 68592 403774 68604
rect 579614 68592 579620 68604
rect 403768 68564 579620 68592
rect 403768 68552 403774 68564
rect 579614 68552 579620 68564
rect 579672 68552 579678 68604
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 35158 68484 35164 68536
rect 35216 68524 35222 68536
rect 87138 68524 87144 68536
rect 35216 68496 87144 68524
rect 35216 68484 35222 68496
rect 87138 68484 87144 68496
rect 87196 68484 87202 68536
<<<<<<< HEAD
rect 193950 68484 193956 68536
rect 194008 68524 194014 68536
rect 430574 68524 430580 68536
rect 194008 68496 430580 68524
rect 194008 68484 194014 68496
rect 430574 68484 430580 68496
rect 430632 68484 430638 68536
=======
rect 177298 68484 177304 68536
rect 177356 68524 177362 68536
rect 229554 68524 229560 68536
rect 177356 68496 229560 68524
rect 177356 68484 177362 68496
rect 229554 68484 229560 68496
rect 229612 68484 229618 68536
rect 244366 68484 244372 68536
rect 244424 68524 244430 68536
rect 245562 68524 245568 68536
rect 244424 68496 245568 68524
rect 244424 68484 244430 68496
rect 245562 68484 245568 68496
rect 245620 68484 245626 68536
rect 295978 68484 295984 68536
rect 296036 68524 296042 68536
rect 488534 68524 488540 68536
rect 296036 68496 488540 68524
rect 296036 68484 296042 68496
rect 488534 68484 488540 68496
rect 488592 68484 488598 68536
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 25498 68416 25504 68468
rect 25556 68456 25562 68468
rect 85758 68456 85764 68468
rect 25556 68428 85764 68456
rect 25556 68416 25562 68428
rect 85758 68416 85764 68428
rect 85816 68416 85822 68468
<<<<<<< HEAD
rect 204438 68416 204444 68468
rect 204496 68456 204502 68468
rect 483014 68456 483020 68468
rect 204496 68428 483020 68456
rect 204496 68416 204502 68428
rect 483014 68416 483020 68428
rect 483072 68416 483078 68468
=======
rect 193950 68416 193956 68468
rect 194008 68456 194014 68468
rect 430574 68456 430580 68468
rect 194008 68428 430580 68456
rect 194008 68416 194014 68428
rect 430574 68416 430580 68428
rect 430632 68416 430638 68468
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 22738 68348 22744 68400
rect 22796 68388 22802 68400
rect 85114 68388 85120 68400
rect 22796 68360 85120 68388
rect 22796 68348 22802 68360
rect 85114 68348 85120 68360
rect 85172 68348 85178 68400
<<<<<<< HEAD
rect 213546 68348 213552 68400
rect 213604 68388 213610 68400
rect 500954 68388 500960 68400
rect 213604 68360 500960 68388
rect 213604 68348 213610 68360
rect 500954 68348 500960 68360
rect 501012 68348 501018 68400
=======
rect 204438 68348 204444 68400
rect 204496 68388 204502 68400
rect 483014 68388 483020 68400
rect 204496 68360 483020 68388
rect 204496 68348 204502 68360
rect 483014 68348 483020 68360
rect 483072 68348 483078 68400
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 50982 68280 50988 68332
rect 51040 68320 51046 68332
rect 111794 68320 111800 68332
rect 51040 68292 111800 68320
rect 51040 68280 51046 68292
rect 111794 68280 111800 68292
rect 111852 68280 111858 68332
<<<<<<< HEAD
rect 134518 68280 134524 68332
rect 134576 68320 134582 68332
rect 312538 68320 312544 68332
rect 134576 68292 312544 68320
rect 134576 68280 134582 68292
rect 312538 68280 312544 68292
rect 312596 68280 312602 68332
rect 314746 68280 314752 68332
rect 314804 68320 314810 68332
rect 315298 68320 315304 68332
rect 314804 68292 315304 68320
rect 314804 68280 314810 68292
rect 315298 68280 315304 68292
rect 315356 68280 315362 68332
rect 404262 68280 404268 68332
rect 404320 68320 404326 68332
rect 579614 68320 579620 68332
rect 404320 68292 579620 68320
rect 404320 68280 404326 68292
rect 579614 68280 579620 68292
rect 579672 68280 579678 68332
=======
rect 213638 68280 213644 68332
rect 213696 68320 213702 68332
rect 500954 68320 500960 68332
rect 213696 68292 500960 68320
rect 213696 68280 213702 68292
rect 500954 68280 500960 68292
rect 501012 68280 501018 68332
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 274358 67260 274364 67312
rect 274416 67300 274422 67312
rect 373994 67300 374000 67312
rect 274416 67272 374000 67300
rect 274416 67260 274422 67272
rect 373994 67260 374000 67272
rect 374052 67260 374058 67312
rect 385126 67260 385132 67312
rect 385184 67300 385190 67312
rect 496814 67300 496820 67312
rect 385184 67272 496820 67300
rect 385184 67260 385190 67272
rect 496814 67260 496820 67272
rect 496872 67260 496878 67312
rect 209038 67192 209044 67244
rect 209096 67232 209102 67244
rect 326522 67232 326528 67244
rect 209096 67204 326528 67232
rect 209096 67192 209102 67204
rect 326522 67192 326528 67204
rect 326580 67192 326586 67244
rect 387242 67192 387248 67244
rect 387300 67232 387306 67244
rect 506474 67232 506480 67244
rect 387300 67204 506480 67232
rect 387300 67192 387306 67204
rect 506474 67192 506480 67204
rect 506532 67192 506538 67244
rect 310146 67124 310152 67176
rect 310204 67164 310210 67176
rect 484394 67164 484400 67176
rect 310204 67136 484400 67164
rect 310204 67124 310210 67136
rect 484394 67124 484400 67136
rect 484452 67124 484458 67176
rect 43438 67056 43444 67108
rect 43496 67096 43502 67108
rect 89806 67096 89812 67108
rect 43496 67068 89812 67096
rect 43496 67056 43502 67068
rect 89806 67056 89812 67068
rect 89864 67056 89870 67108
rect 292390 67056 292396 67108
rect 292448 67096 292454 67108
rect 466454 67096 466460 67108
rect 292448 67068 466460 67096
rect 292448 67056 292454 67068
rect 466454 67056 466460 67068
rect 466512 67056 466518 67108
rect 39298 66988 39304 67040
rect 39356 67028 39362 67040
rect 88518 67028 88524 67040
rect 39356 67000 88524 67028
rect 39356 66988 39362 67000
rect 88518 66988 88524 67000
rect 88576 66988 88582 67040
rect 192570 66988 192576 67040
rect 192628 67028 192634 67040
rect 423674 67028 423680 67040
rect 192628 67000 423680 67028
rect 192628 66988 192634 67000
rect 423674 66988 423680 67000
rect 423732 66988 423738 67040
rect 32398 66920 32404 66972
rect 32456 66960 32462 66972
rect 86494 66960 86500 66972
rect 32456 66932 86500 66960
rect 32456 66920 32462 66932
rect 86494 66920 86500 66932
rect 86552 66920 86558 66972
rect 205818 66920 205824 66972
rect 205876 66960 205882 66972
rect 489914 66960 489920 66972
rect 205876 66932 489920 66960
rect 205876 66920 205882 66932
rect 489914 66920 489920 66932
rect 489972 66920 489978 66972
rect 15838 66852 15844 66904
rect 15896 66892 15902 66904
rect 107378 66892 107384 66904
rect 15896 66864 107384 66892
rect 15896 66852 15902 66864
rect 107378 66852 107384 66864
rect 107436 66852 107442 66904
rect 209314 66852 209320 66904
rect 209372 66892 209378 66904
rect 507854 66892 507860 66904
rect 209372 66864 507860 66892
rect 209372 66852 209378 66864
rect 507854 66852 507860 66864
rect 507912 66852 507918 66904
rect 387978 65832 387984 65884
rect 388036 65872 388042 65884
rect 510614 65872 510620 65884
rect 388036 65844 510620 65872
rect 388036 65832 388042 65844
rect 510614 65832 510620 65844
rect 510672 65832 510678 65884
<<<<<<< HEAD
rect 392394 65764 392400 65816
rect 392452 65804 392458 65816
rect 524414 65804 524420 65816
rect 392452 65776 524420 65804
rect 392452 65764 392458 65776
=======
rect 391934 65764 391940 65816
rect 391992 65804 391998 65816
rect 524414 65804 524420 65816
rect 391992 65776 524420 65804
rect 391992 65764 391998 65776
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 524414 65764 524420 65776
rect 524472 65764 524478 65816
rect 289538 65696 289544 65748
rect 289596 65736 289602 65748
rect 463694 65736 463700 65748
rect 289596 65708 463700 65736
rect 289596 65696 289602 65708
rect 463694 65696 463700 65708
rect 463752 65696 463758 65748
rect 82354 65628 82360 65680
rect 82412 65668 82418 65680
rect 114646 65668 114652 65680
rect 82412 65640 114652 65668
rect 82412 65628 82418 65640
rect 114646 65628 114652 65640
rect 114704 65628 114710 65680
rect 293770 65628 293776 65680
rect 293828 65668 293834 65680
rect 470594 65668 470600 65680
rect 293828 65640 470600 65668
rect 293828 65628 293834 65640
rect 470594 65628 470600 65640
rect 470652 65628 470658 65680
rect 197446 65560 197452 65612
rect 197504 65600 197510 65612
rect 448514 65600 448520 65612
rect 197504 65572 448520 65600
rect 197504 65560 197510 65572
rect 448514 65560 448520 65572
rect 448572 65560 448578 65612
rect 53650 65492 53656 65544
rect 53708 65532 53714 65544
rect 115106 65532 115112 65544
rect 53708 65504 115112 65532
rect 53708 65492 53714 65504
rect 115106 65492 115112 65504
rect 115164 65492 115170 65544
rect 222562 65492 222568 65544
rect 222620 65532 222626 65544
rect 575474 65532 575480 65544
rect 222620 65504 575480 65532
rect 222620 65492 222626 65504
rect 575474 65492 575480 65504
rect 575532 65492 575538 65544
rect 383470 64336 383476 64388
rect 383528 64376 383534 64388
rect 485774 64376 485780 64388
rect 383528 64348 485780 64376
rect 383528 64336 383534 64348
rect 485774 64336 485780 64348
rect 485832 64336 485838 64388
rect 390370 64268 390376 64320
rect 390428 64308 390434 64320
rect 517514 64308 517520 64320
rect 390428 64280 517520 64308
rect 390428 64268 390434 64280
rect 517514 64268 517520 64280
rect 517572 64268 517578 64320
rect 394510 64200 394516 64252
rect 394568 64240 394574 64252
rect 539594 64240 539600 64252
rect 394568 64212 539600 64240
rect 394568 64200 394574 64212
rect 539594 64200 539600 64212
rect 539652 64200 539658 64252
rect 288250 64132 288256 64184
rect 288308 64172 288314 64184
rect 456886 64172 456892 64184
rect 288308 64144 456892 64172
rect 288308 64132 288314 64144
rect 456886 64132 456892 64144
rect 456944 64132 456950 64184
rect 393130 62840 393136 62892
rect 393188 62880 393194 62892
rect 530578 62880 530584 62892
rect 393188 62852 530584 62880
rect 393188 62840 393194 62852
rect 530578 62840 530584 62852
rect 530636 62840 530642 62892
rect 395890 62772 395896 62824
rect 395948 62812 395954 62824
rect 546494 62812 546500 62824
rect 395948 62784 546500 62812
rect 395948 62772 395954 62784
rect 546494 62772 546500 62784
rect 546552 62772 546558 62824
rect 406746 60664 406752 60716
rect 406804 60704 406810 60716
rect 580166 60704 580172 60716
rect 406804 60676 580172 60704
rect 406804 60664 406810 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 389082 58624 389088 58676
rect 389140 58664 389146 58676
rect 514754 58664 514760 58676
rect 389140 58636 514760 58664
rect 389140 58624 389146 58636
rect 514754 58624 514760 58636
rect 514812 58624 514818 58676
rect 235902 50328 235908 50380
rect 235960 50368 235966 50380
rect 331858 50368 331864 50380
rect 235960 50340 331864 50368
rect 235960 50328 235966 50340
rect 331858 50328 331864 50340
rect 331916 50328 331922 50380
rect 394602 50328 394608 50380
rect 394660 50368 394666 50380
rect 542354 50368 542360 50380
rect 394660 50340 542360 50368
rect 394660 50328 394666 50340
rect 542354 50328 542360 50340
rect 542412 50328 542418 50380
rect 45370 48968 45376 49020
rect 45428 49008 45434 49020
rect 87598 49008 87604 49020
rect 45428 48980 87604 49008
rect 45428 48968 45434 48980
rect 87598 48968 87604 48980
rect 87656 48968 87662 49020
rect 176470 48968 176476 49020
rect 176528 49008 176534 49020
rect 338298 49008 338304 49020
rect 176528 48980 338304 49008
rect 176528 48968 176534 48980
rect 338298 48968 338304 48980
rect 338356 48968 338362 49020
rect 175090 47540 175096 47592
rect 175148 47580 175154 47592
rect 331306 47580 331312 47592
rect 175148 47552 331312 47580
rect 175148 47540 175154 47552
rect 331306 47540 331312 47552
rect 331364 47540 331370 47592
rect 406654 46860 406660 46912
rect 406712 46900 406718 46912
rect 580166 46900 580172 46912
rect 406712 46872 580172 46900
rect 406712 46860 406718 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 228450 44820 228456 44872
rect 228508 44860 228514 44872
rect 328546 44860 328552 44872
rect 228508 44832 328552 44860
rect 228508 44820 228514 44832
rect 328546 44820 328552 44832
rect 328604 44820 328610 44872
rect 406562 33056 406568 33108
rect 406620 33096 406626 33108
rect 579890 33096 579896 33108
rect 406620 33068 579896 33096
rect 406620 33056 406626 33068
rect 579890 33056 579896 33068
rect 579948 33056 579954 33108
rect 238018 25508 238024 25560
rect 238076 25548 238082 25560
rect 331398 25548 331404 25560
rect 238076 25520 331404 25548
rect 238076 25508 238082 25520
rect 331398 25508 331404 25520
rect 331456 25508 331462 25560
rect 289722 24080 289728 24132
rect 289780 24120 289786 24132
rect 459554 24120 459560 24132
rect 289780 24092 459560 24120
rect 289780 24080 289786 24092
rect 459554 24080 459560 24092
rect 459612 24080 459618 24132
rect 227070 22720 227076 22772
rect 227128 22760 227134 22772
rect 329926 22760 329932 22772
rect 227128 22732 329932 22760
rect 227128 22720 227134 22732
rect 329926 22720 329932 22732
rect 329984 22720 329990 22772
rect 393222 22720 393228 22772
rect 393280 22760 393286 22772
rect 535454 22760 535460 22772
rect 393280 22732 535460 22760
rect 393280 22720 393286 22732
rect 535454 22720 535460 22732
rect 535512 22720 535518 22772
rect 268930 21360 268936 21412
rect 268988 21400 268994 21412
rect 354030 21400 354036 21412
rect 268988 21372 354036 21400
rect 268988 21360 268994 21372
rect 354030 21360 354036 21372
rect 354088 21360 354094 21412
rect 390462 21360 390468 21412
rect 390520 21400 390526 21412
rect 521654 21400 521660 21412
rect 390520 21372 521660 21400
rect 390520 21360 390526 21372
rect 521654 21360 521660 21372
rect 521712 21360 521718 21412
rect 406470 20612 406476 20664
rect 406528 20652 406534 20664
rect 579890 20652 579896 20664
rect 406528 20624 579896 20652
rect 406528 20612 406534 20624
rect 579890 20612 579896 20624
rect 579948 20612 579954 20664
rect 295978 19932 295984 19984
rect 296036 19972 296042 19984
rect 342346 19972 342352 19984
rect 296036 19944 342352 19972
rect 296036 19932 296042 19944
rect 342346 19932 342352 19944
rect 342404 19932 342410 19984
rect 198550 18776 198556 18828
rect 198608 18816 198614 18828
rect 236086 18816 236092 18828
rect 198608 18788 236092 18816
rect 198608 18776 198614 18788
rect 236086 18776 236092 18788
rect 236144 18776 236150 18828
rect 222930 18708 222936 18760
rect 222988 18748 222994 18760
rect 329834 18748 329840 18760
rect 222988 18720 329840 18748
rect 222988 18708 222994 18720
rect 329834 18708 329840 18720
rect 329892 18708 329898 18760
rect 202598 18640 202604 18692
rect 202656 18680 202662 18692
rect 327166 18680 327172 18692
rect 202656 18652 327172 18680
rect 202656 18640 202662 18652
rect 327166 18640 327172 18652
rect 327224 18640 327230 18692
rect 162118 18572 162124 18624
rect 162176 18612 162182 18624
rect 313274 18612 313280 18624
rect 162176 18584 313280 18612
rect 162176 18572 162182 18584
rect 313274 18572 313280 18584
rect 313332 18572 313338 18624
rect 386322 18572 386328 18624
rect 386380 18612 386386 18624
rect 499574 18612 499580 18624
rect 386380 18584 499580 18612
rect 386380 18572 386386 18584
rect 499574 18572 499580 18584
rect 499632 18572 499638 18624
rect 249058 17892 249064 17944
rect 249116 17932 249122 17944
rect 251174 17932 251180 17944
rect 249116 17904 251180 17932
rect 249116 17892 249122 17904
rect 251174 17892 251180 17904
rect 251232 17892 251238 17944
rect 242250 17552 242256 17604
rect 242308 17592 242314 17604
rect 334066 17592 334072 17604
rect 242308 17564 334072 17592
rect 242308 17552 242314 17564
rect 334066 17552 334072 17564
rect 334124 17552 334130 17604
rect 271690 17484 271696 17536
rect 271748 17524 271754 17536
rect 367094 17524 367100 17536
rect 271748 17496 367100 17524
rect 271748 17484 271754 17496
rect 367094 17484 367100 17496
rect 367152 17484 367158 17536
rect 177850 17416 177856 17468
rect 177908 17456 177914 17468
rect 231946 17456 231952 17468
rect 177908 17428 231952 17456
rect 177908 17416 177914 17428
rect 231946 17416 231952 17428
rect 232004 17416 232010 17468
rect 232590 17416 232596 17468
rect 232648 17456 232654 17468
rect 328454 17456 328460 17468
rect 232648 17428 328460 17456
rect 232648 17416 232654 17428
rect 328454 17416 328460 17428
rect 328512 17416 328518 17468
rect 195238 17348 195244 17400
rect 195296 17388 195302 17400
rect 324406 17388 324412 17400
rect 195296 17360 324412 17388
rect 195296 17348 195302 17360
rect 324406 17348 324412 17360
rect 324464 17348 324470 17400
rect 178678 17280 178684 17332
rect 178736 17320 178742 17332
rect 320358 17320 320364 17332
rect 178736 17292 320364 17320
rect 178736 17280 178742 17292
rect 320358 17280 320364 17292
rect 320416 17280 320422 17332
rect 175090 17212 175096 17264
rect 175148 17252 175154 17264
rect 321646 17252 321652 17264
rect 175148 17224 321652 17252
rect 175148 17212 175154 17224
rect 321646 17212 321652 17224
rect 321704 17212 321710 17264
rect 383562 17212 383568 17264
rect 383620 17252 383626 17264
rect 481726 17252 481732 17264
rect 383620 17224 481732 17252
rect 383620 17212 383626 17224
rect 481726 17212 481732 17224
rect 481784 17212 481790 17264
rect 270310 16328 270316 16380
rect 270368 16368 270374 16380
rect 354122 16368 354128 16380
rect 270368 16340 354128 16368
rect 270368 16328 270374 16340
rect 354122 16328 354128 16340
rect 354180 16328 354186 16380
rect 271782 16260 271788 16312
rect 271840 16300 271846 16312
<<<<<<< HEAD
rect 371694 16300 371700 16312
rect 271840 16272 371700 16300
rect 271840 16260 271846 16272
rect 371694 16260 371700 16272
rect 371752 16260 371758 16312
=======
rect 371234 16300 371240 16312
rect 271840 16272 371240 16300
rect 271840 16260 271846 16272
rect 371234 16260 371240 16272
rect 371292 16260 371298 16312
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 224402 16192 224408 16244
rect 224460 16232 224466 16244
rect 327074 16232 327080 16244
rect 224460 16204 327080 16232
rect 224460 16192 224466 16204
rect 327074 16192 327080 16204
rect 327132 16192 327138 16244
rect 196618 16124 196624 16176
rect 196676 16164 196682 16176
rect 323118 16164 323124 16176
rect 196676 16136 323124 16164
rect 196676 16124 196682 16136
rect 323118 16124 323124 16136
rect 323176 16124 323182 16176
rect 173250 16056 173256 16108
rect 173308 16096 173314 16108
rect 313458 16096 313464 16108
rect 173308 16068 313464 16096
rect 173308 16056 173314 16068
rect 313458 16056 313464 16068
rect 313516 16056 313522 16108
rect 173158 15988 173164 16040
rect 173216 16028 173222 16040
rect 316310 16028 316316 16040
rect 173216 16000 316316 16028
rect 173216 15988 173222 16000
rect 316310 15988 316316 16000
rect 316368 15988 316374 16040
rect 164142 15920 164148 15972
rect 164200 15960 164206 15972
rect 309778 15960 309784 15972
rect 164200 15932 309784 15960
rect 164200 15920 164206 15932
rect 309778 15920 309784 15932
rect 309836 15920 309842 15972
rect 197170 15852 197176 15904
rect 197228 15892 197234 15904
rect 441522 15892 441528 15904
rect 197228 15864 441528 15892
rect 197228 15852 197234 15864
rect 441522 15852 441528 15864
rect 441580 15852 441586 15904
rect 267550 14968 267556 15020
rect 267608 15008 267614 15020
rect 349338 15008 349344 15020
rect 267608 14980 349344 15008
rect 267608 14968 267614 14980
rect 349338 14968 349344 14980
rect 349396 14968 349402 15020
rect 231210 14900 231216 14952
rect 231268 14940 231274 14952
rect 331214 14940 331220 14952
rect 231268 14912 331220 14940
rect 231268 14900 231274 14912
rect 331214 14900 331220 14912
rect 331272 14900 331278 14952
rect 206370 14832 206376 14884
rect 206428 14872 206434 14884
rect 324314 14872 324320 14884
rect 206428 14844 324320 14872
rect 206428 14832 206434 14844
rect 324314 14832 324320 14844
rect 324372 14832 324378 14884
rect 195330 14764 195336 14816
rect 195388 14804 195394 14816
rect 321554 14804 321560 14816
rect 195388 14776 321560 14804
rect 195388 14764 195394 14776
rect 321554 14764 321560 14776
rect 321612 14764 321618 14816
rect 170950 14696 170956 14748
rect 171008 14736 171014 14748
<<<<<<< HEAD
rect 310238 14736 310244 14748
rect 171008 14708 310244 14736
rect 171008 14696 171014 14708
rect 310238 14696 310244 14708
rect 310296 14696 310302 14748
rect 175182 14628 175188 14680
rect 175240 14668 175246 14680
rect 335078 14668 335084 14680
rect 175240 14640 335084 14668
rect 175240 14628 175246 14640
rect 335078 14628 335084 14640
rect 335136 14628 335142 14680
=======
rect 309778 14736 309784 14748
rect 171008 14708 309784 14736
rect 171008 14696 171014 14708
rect 309778 14696 309784 14708
rect 309836 14696 309842 14748
rect 175182 14628 175188 14680
rect 175240 14668 175246 14680
rect 334618 14668 334624 14680
rect 175240 14640 334624 14668
rect 175240 14628 175246 14640
rect 334618 14628 334624 14640
rect 334676 14628 334682 14680
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 179230 14560 179236 14612
rect 179288 14600 179294 14612
rect 352834 14600 352840 14612
rect 179288 14572 352840 14600
rect 179288 14560 179294 14572
rect 352834 14560 352840 14572
rect 352892 14560 352898 14612
rect 170398 14492 170404 14544
rect 170456 14532 170462 14544
rect 230566 14532 230572 14544
rect 170456 14504 230572 14532
rect 170456 14492 170462 14504
rect 230566 14492 230572 14504
rect 230624 14492 230630 14544
rect 292482 14492 292488 14544
rect 292540 14532 292546 14544
rect 478138 14532 478144 14544
rect 292540 14504 478144 14532
rect 292540 14492 292546 14504
rect 478138 14492 478144 14504
rect 478196 14492 478202 14544
rect 30098 14424 30104 14476
rect 30156 14464 30162 14476
rect 64966 14464 64972 14476
rect 30156 14436 64972 14464
rect 30156 14424 30162 14436
rect 64966 14424 64972 14436
rect 65024 14424 65030 14476
rect 195790 14424 195796 14476
rect 195848 14464 195854 14476
<<<<<<< HEAD
rect 437934 14464 437940 14476
rect 195848 14436 437940 14464
rect 195848 14424 195854 14436
rect 437934 14424 437940 14436
rect 437992 14424 437998 14476
=======
rect 437474 14464 437480 14476
rect 195848 14436 437480 14464
rect 195848 14424 195854 14436
rect 437474 14424 437480 14436
rect 437532 14424 437538 14476
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 104158 14084 104164 14136
rect 104216 14124 104222 14136
rect 105722 14124 105728 14136
rect 104216 14096 105728 14124
rect 104216 14084 104222 14096
rect 105722 14084 105728 14096
rect 105780 14084 105786 14136
rect 173618 13676 173624 13728
rect 173676 13716 173682 13728
rect 231854 13716 231860 13728
rect 173676 13688 231860 13716
rect 173676 13676 173682 13688
rect 231854 13676 231860 13688
rect 231912 13676 231918 13728
rect 270402 13676 270408 13728
rect 270460 13716 270466 13728
rect 360838 13716 360844 13728
rect 270460 13688 360844 13716
rect 270460 13676 270466 13688
rect 360838 13676 360844 13688
rect 360896 13676 360902 13728
rect 195606 13608 195612 13660
rect 195664 13648 195670 13660
rect 287698 13648 287704 13660
rect 195664 13620 287704 13648
rect 195664 13608 195670 13620
rect 287698 13608 287704 13620
rect 287756 13608 287762 13660
rect 231762 13540 231768 13592
rect 231820 13580 231826 13592
rect 327718 13580 327724 13592
rect 231820 13552 327724 13580
rect 231820 13540 231826 13552
rect 327718 13540 327724 13552
rect 327776 13540 327782 13592
rect 169570 13472 169576 13524
rect 169628 13512 169634 13524
<<<<<<< HEAD
rect 306742 13512 306748 13524
rect 169628 13484 306748 13512
rect 169628 13472 169634 13484
rect 306742 13472 306748 13484
rect 306800 13472 306806 13524
=======
rect 306374 13512 306380 13524
rect 169628 13484 306380 13512
rect 169628 13472 169634 13484
rect 306374 13472 306380 13484
rect 306432 13472 306438 13524
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 173802 13404 173808 13456
rect 173860 13444 173866 13456
rect 324406 13444 324412 13456
rect 173860 13416 324412 13444
rect 173860 13404 173866 13416
rect 324406 13404 324412 13416
rect 324464 13404 324470 13456
rect 173710 13336 173716 13388
rect 173768 13376 173774 13388
rect 327994 13376 328000 13388
rect 173768 13348 328000 13376
rect 173768 13336 173774 13348
rect 327994 13336 328000 13348
rect 328052 13336 328058 13388
rect 177758 13268 177764 13320
rect 177816 13308 177822 13320
rect 349246 13308 349252 13320
rect 177816 13280 349252 13308
rect 177816 13268 177822 13280
rect 349246 13268 349252 13280
rect 349304 13268 349310 13320
rect 195882 13200 195888 13252
rect 195940 13240 195946 13252
<<<<<<< HEAD
rect 434438 13240 434444 13252
rect 195940 13212 434444 13240
rect 195940 13200 195946 13212
rect 434438 13200 434444 13212
rect 434496 13200 434502 13252
rect 198642 13132 198648 13184
rect 198700 13172 198706 13184
rect 452102 13172 452108 13184
rect 198700 13144 452108 13172
rect 198700 13132 198706 13144
rect 452102 13132 452108 13144
rect 452160 13132 452166 13184
=======
rect 433978 13240 433984 13252
rect 195940 13212 433984 13240
rect 195940 13200 195946 13212
rect 433978 13200 433984 13212
rect 434036 13200 434042 13252
rect 198642 13132 198648 13184
rect 198700 13172 198706 13184
rect 451642 13172 451648 13184
rect 198700 13144 451648 13172
rect 198700 13132 198706 13144
rect 451642 13132 451648 13144
rect 451700 13132 451706 13184
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 206922 13064 206928 13116
rect 206980 13104 206986 13116
rect 494698 13104 494704 13116
rect 206980 13076 494704 13104
rect 206980 13064 206986 13076
rect 494698 13064 494704 13076
rect 494756 13064 494762 13116
rect 267642 12384 267648 12436
rect 267700 12424 267706 12436
rect 346946 12424 346952 12436
rect 267700 12396 346952 12424
rect 267700 12384 267706 12396
rect 346946 12384 346952 12396
rect 347004 12384 347010 12436
rect 181898 12316 181904 12368
rect 181956 12356 181962 12368
rect 291838 12356 291844 12368
rect 181956 12328 291844 12356
rect 181956 12316 181962 12328
rect 291838 12316 291844 12328
rect 291896 12316 291902 12368
rect 169662 12248 169668 12300
rect 169720 12288 169726 12300
rect 303154 12288 303160 12300
rect 169720 12260 303160 12288
rect 169720 12248 169726 12260
rect 303154 12248 303160 12260
rect 303212 12248 303218 12300
rect 171042 12180 171048 12232
rect 171100 12220 171106 12232
rect 313826 12220 313832 12232
rect 171100 12192 313832 12220
rect 171100 12180 171106 12192
rect 313826 12180 313832 12192
rect 313884 12180 313890 12232
rect 169570 12112 169576 12164
rect 169628 12152 169634 12164
rect 230474 12152 230480 12164
rect 169628 12124 230480 12152
rect 169628 12112 169634 12124
rect 230474 12112 230480 12124
rect 230532 12112 230538 12164
rect 286870 12112 286876 12164
rect 286928 12152 286934 12164
<<<<<<< HEAD
rect 446214 12152 446220 12164
rect 286928 12124 446220 12152
rect 286928 12112 286934 12124
rect 446214 12112 446220 12124
rect 446272 12112 446278 12164
=======
rect 445754 12152 445760 12164
rect 286928 12124 445760 12152
rect 286928 12112 286934 12124
rect 445754 12112 445760 12124
rect 445812 12112 445818 12164
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 160738 12044 160744 12096
rect 160796 12084 160802 12096
rect 227806 12084 227812 12096
rect 160796 12056 227812 12084
rect 160796 12044 160802 12056
rect 227806 12044 227812 12056
rect 227864 12044 227870 12096
rect 286962 12044 286968 12096
rect 287020 12084 287026 12096
rect 449802 12084 449808 12096
rect 287020 12056 449808 12084
rect 287020 12044 287026 12056
rect 449802 12044 449808 12056
rect 449860 12044 449866 12096
rect 162670 11976 162676 12028
rect 162728 12016 162734 12028
rect 267734 12016 267740 12028
rect 162728 11988 267740 12016
rect 162728 11976 162734 11988
rect 267734 11976 267740 11988
rect 267792 11976 267798 12028
rect 288342 11976 288348 12028
rect 288400 12016 288406 12028
rect 453298 12016 453304 12028
rect 288400 11988 453304 12016
rect 288400 11976 288406 11988
rect 453298 11976 453304 11988
rect 453356 11976 453362 12028
rect 176562 11908 176568 11960
rect 176620 11948 176626 11960
rect 341058 11948 341064 11960
rect 176620 11920 341064 11948
rect 176620 11908 176626 11920
rect 341058 11908 341064 11920
rect 341116 11908 341122 11960
rect 353938 11908 353944 11960
rect 353996 11948 354002 11960
<<<<<<< HEAD
rect 427262 11948 427268 11960
rect 353996 11920 427268 11948
rect 353996 11908 354002 11920
rect 427262 11908 427268 11920
rect 427320 11908 427326 11960
rect 165522 11840 165528 11892
rect 165580 11880 165586 11892
rect 285398 11880 285404 11892
rect 165580 11852 285404 11880
rect 165580 11840 165586 11852
rect 285398 11840 285404 11852
rect 285456 11840 285462 11892
rect 296622 11840 296628 11892
rect 296680 11880 296686 11892
rect 499390 11880 499396 11892
rect 296680 11852 499396 11880
rect 296680 11840 296686 11852
rect 499390 11840 499396 11852
rect 499448 11840 499454 11892
=======
rect 426802 11948 426808 11960
rect 353996 11920 426808 11948
rect 353996 11908 354002 11920
rect 426802 11908 426808 11920
rect 426860 11908 426866 11960
rect 165522 11840 165528 11892
rect 165580 11880 165586 11892
rect 284938 11880 284944 11892
rect 165580 11852 284944 11880
rect 165580 11840 165586 11852
rect 284938 11840 284944 11852
rect 284996 11840 285002 11892
rect 296622 11840 296628 11892
rect 296680 11880 296686 11892
rect 498930 11880 498936 11892
rect 296680 11852 498936 11880
rect 296680 11840 296686 11852
rect 498930 11840 498936 11852
rect 498988 11840 498994 11892
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 197262 11772 197268 11824
rect 197320 11812 197326 11824
rect 445018 11812 445024 11824
rect 197320 11784 445024 11812
rect 197320 11772 197326 11784
rect 445018 11772 445024 11784
rect 445076 11772 445082 11824
rect 224310 11704 224316 11756
rect 224368 11744 224374 11756
rect 498194 11744 498200 11756
rect 224368 11716 498200 11744
rect 224368 11704 224374 11716
rect 498194 11704 498200 11716
rect 498252 11704 498258 11756
rect 226978 11636 226984 11688
rect 227036 11676 227042 11688
<<<<<<< HEAD
rect 281902 11676 281908 11688
rect 227036 11648 281908 11676
rect 227036 11636 227042 11648
rect 281902 11636 281908 11648
rect 281960 11636 281966 11688
=======
rect 281534 11676 281540 11688
rect 227036 11648 281540 11676
rect 227036 11636 227042 11648
rect 281534 11636 281540 11648
rect 281592 11636 281598 11688
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 278682 10956 278688 11008
rect 278740 10996 278746 11008
rect 407206 10996 407212 11008
rect 278740 10968 407212 10996
rect 278740 10956 278746 10968
rect 407206 10956 407212 10968
rect 407264 10956 407270 11008
rect 202506 10888 202512 10940
rect 202564 10928 202570 10940
rect 237466 10928 237472 10940
rect 202564 10900 237472 10928
rect 202564 10888 202570 10900
rect 237466 10888 237472 10900
rect 237524 10888 237530 10940
rect 279970 10888 279976 10940
rect 280028 10928 280034 10940
rect 410794 10928 410800 10940
rect 280028 10900 410800 10928
rect 280028 10888 280034 10900
rect 410794 10888 410800 10900
rect 410852 10888 410858 10940
rect 191558 10820 191564 10872
rect 191616 10860 191622 10872
rect 234706 10860 234712 10872
rect 191616 10832 234712 10860
rect 191616 10820 191622 10832
rect 234706 10820 234712 10832
rect 234764 10820 234770 10872
rect 280062 10820 280068 10872
rect 280120 10860 280126 10872
rect 414290 10860 414296 10872
rect 280120 10832 414296 10860
rect 280120 10820 280126 10832
rect 414290 10820 414296 10832
rect 414348 10820 414354 10872
rect 414658 10820 414664 10872
rect 414716 10860 414722 10872
rect 490006 10860 490012 10872
rect 414716 10832 490012 10860
rect 414716 10820 414722 10832
rect 490006 10820 490012 10832
rect 490064 10820 490070 10872
rect 187326 10752 187332 10804
rect 187384 10792 187390 10804
rect 232498 10792 232504 10804
rect 187384 10764 232504 10792
rect 187384 10752 187390 10764
rect 232498 10752 232504 10764
rect 232556 10752 232562 10804
rect 281350 10752 281356 10804
rect 281408 10792 281414 10804
<<<<<<< HEAD
rect 417878 10792 417884 10804
rect 281408 10764 417884 10792
rect 281408 10752 281414 10764
rect 417878 10752 417884 10764
rect 417936 10752 417942 10804
=======
rect 417418 10792 417424 10804
rect 281408 10764 417424 10792
rect 281408 10752 281414 10764
rect 417418 10752 417424 10764
rect 417476 10752 417482 10804
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 209130 10684 209136 10736
rect 209188 10724 209194 10736
rect 274818 10724 274824 10736
rect 209188 10696 274824 10724
rect 209188 10684 209194 10696
rect 274818 10684 274824 10696
rect 274876 10684 274882 10736
rect 281258 10684 281264 10736
rect 281316 10724 281322 10736
<<<<<<< HEAD
rect 421374 10724 421380 10736
rect 281316 10696 421380 10724
rect 281316 10684 281322 10696
rect 421374 10684 421380 10696
rect 421432 10684 421438 10736
=======
rect 420914 10724 420920 10736
rect 281316 10696 420920 10724
rect 281316 10684 281322 10696
rect 420914 10684 420920 10696
rect 420972 10684 420978 10736
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 162486 10616 162492 10668
rect 162544 10656 162550 10668
rect 228358 10656 228364 10668
rect 162544 10628 228364 10656
rect 162544 10616 162550 10628
rect 228358 10616 228364 10628
rect 228416 10616 228422 10668
rect 282730 10616 282736 10668
rect 282788 10656 282794 10668
rect 424962 10656 424968 10668
rect 282788 10628 424968 10656
rect 282788 10616 282794 10628
rect 424962 10616 424968 10628
rect 425020 10616 425026 10668
rect 158622 10548 158628 10600
rect 158680 10588 158686 10600
rect 249978 10588 249984 10600
rect 158680 10560 249984 10588
rect 158680 10548 158686 10560
rect 249978 10548 249984 10560
rect 250036 10548 250042 10600
rect 250438 10548 250444 10600
rect 250496 10588 250502 10600
rect 278314 10588 278320 10600
rect 250496 10560 278320 10588
rect 250496 10548 250502 10560
rect 278314 10548 278320 10560
rect 278372 10548 278378 10600
rect 282822 10548 282828 10600
rect 282880 10588 282886 10600
rect 428458 10588 428464 10600
rect 282880 10560 428464 10588
rect 282880 10548 282886 10560
rect 428458 10548 428464 10560
rect 428516 10548 428522 10600
rect 159910 10480 159916 10532
rect 159968 10520 159974 10532
rect 253474 10520 253480 10532
rect 159968 10492 253480 10520
rect 159968 10480 159974 10492
rect 253474 10480 253480 10492
rect 253532 10480 253538 10532
rect 284202 10480 284208 10532
rect 284260 10520 284266 10532
rect 432046 10520 432052 10532
rect 284260 10492 432052 10520
rect 284260 10480 284266 10492
rect 432046 10480 432052 10492
rect 432104 10480 432110 10532
rect 161382 10412 161388 10464
rect 161440 10452 161446 10464
<<<<<<< HEAD
rect 259454 10452 259460 10464
rect 161440 10424 259460 10452
rect 161440 10412 161446 10424
rect 259454 10412 259460 10424
rect 259512 10412 259518 10464
rect 284110 10412 284116 10464
rect 284168 10452 284174 10464
rect 435542 10452 435548 10464
rect 284168 10424 435548 10452
rect 284168 10412 284174 10424
rect 435542 10412 435548 10424
rect 435600 10412 435606 10464
=======
rect 260650 10452 260656 10464
rect 161440 10424 260656 10452
rect 161440 10412 161446 10424
rect 260650 10412 260656 10424
rect 260708 10412 260714 10464
rect 284110 10412 284116 10464
rect 284168 10452 284174 10464
rect 435082 10452 435088 10464
rect 284168 10424 435088 10452
rect 284168 10412 284174 10424
rect 435082 10412 435088 10424
rect 435140 10412 435146 10464
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 161290 10344 161296 10396
rect 161348 10384 161354 10396
rect 264146 10384 264152 10396
rect 161348 10356 264152 10384
rect 161348 10344 161354 10356
rect 264146 10344 264152 10356
rect 264204 10344 264210 10396
rect 285490 10344 285496 10396
rect 285548 10384 285554 10396
rect 439130 10384 439136 10396
rect 285548 10356 439136 10384
rect 285548 10344 285554 10356
rect 439130 10344 439136 10356
rect 439188 10344 439194 10396
rect 162762 10276 162768 10328
rect 162820 10316 162826 10328
<<<<<<< HEAD
rect 271230 10316 271236 10328
rect 162820 10288 271236 10316
rect 162820 10276 162826 10288
rect 271230 10276 271236 10288
rect 271288 10276 271294 10328
=======
rect 270770 10316 270776 10328
rect 162820 10288 270776 10316
rect 162820 10276 162826 10288
rect 270770 10276 270776 10288
rect 270828 10276 270834 10328
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 285582 10276 285588 10328
rect 285640 10316 285646 10328
rect 442626 10316 442632 10328
rect 285640 10288 442632 10316
rect 285640 10276 285646 10288
rect 442626 10276 442632 10288
rect 442684 10276 442690 10328
rect 278590 10208 278596 10260
rect 278648 10248 278654 10260
rect 403618 10248 403624 10260
rect 278648 10220 403624 10248
rect 278648 10208 278654 10220
rect 403618 10208 403624 10220
rect 403676 10208 403682 10260
rect 277302 10140 277308 10192
rect 277360 10180 277366 10192
rect 398834 10180 398840 10192
rect 277360 10152 398840 10180
rect 277360 10140 277366 10152
rect 398834 10140 398840 10152
rect 398892 10140 398898 10192
rect 277210 10072 277216 10124
rect 277268 10112 277274 10124
<<<<<<< HEAD
rect 396534 10112 396540 10124
rect 277268 10084 396540 10112
rect 277268 10072 277274 10084
rect 396534 10072 396540 10084
rect 396592 10072 396598 10124
rect 275922 10004 275928 10056
rect 275980 10044 275986 10056
rect 393038 10044 393044 10056
rect 275980 10016 393044 10044
rect 275980 10004 275986 10016
rect 393038 10004 393044 10016
rect 393096 10004 393102 10056
=======
rect 396074 10112 396080 10124
rect 277268 10084 396080 10112
rect 277268 10072 277274 10084
rect 396074 10072 396080 10084
rect 396132 10072 396138 10124
rect 275922 10004 275928 10056
rect 275980 10044 275986 10056
rect 392578 10044 392584 10056
rect 275980 10016 392584 10044
rect 275980 10004 275986 10016
rect 392578 10004 392584 10016
rect 392636 10004 392642 10056
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 275830 9936 275836 9988
rect 275888 9976 275894 9988
rect 389450 9976 389456 9988
rect 275888 9948 389456 9976
rect 275888 9936 275894 9948
rect 389450 9936 389456 9948
rect 389508 9936 389514 9988
rect 274542 9868 274548 9920
rect 274600 9908 274606 9920
rect 385954 9908 385960 9920
rect 274600 9880 385960 9908
rect 274600 9868 274606 9880
rect 385954 9868 385960 9880
rect 386012 9868 386018 9920
rect 274450 9800 274456 9852
rect 274508 9840 274514 9852
rect 382366 9840 382372 9852
rect 274508 9812 382372 9840
rect 274508 9800 274514 9812
rect 382366 9800 382372 9812
rect 382424 9800 382430 9852
rect 273162 9732 273168 9784
rect 273220 9772 273226 9784
<<<<<<< HEAD
rect 378870 9772 378876 9784
rect 273220 9744 378876 9772
rect 273220 9732 273226 9744
rect 378870 9732 378876 9744
rect 378928 9732 378934 9784
=======
rect 378410 9772 378416 9784
rect 273220 9744 378416 9772
rect 273220 9732 273226 9744
rect 378410 9732 378416 9744
rect 378468 9732 378474 9784
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 215662 9596 215668 9648
rect 215720 9636 215726 9648
rect 240226 9636 240232 9648
rect 215720 9608 240232 9636
rect 215720 9596 215726 9608
rect 240226 9596 240232 9608
rect 240284 9596 240290 9648
rect 240502 9596 240508 9648
rect 240560 9636 240566 9648
rect 244366 9636 244372 9648
rect 240560 9608 244372 9636
rect 240560 9596 240566 9608
rect 244366 9596 244372 9608
rect 244424 9596 244430 9648
rect 308950 9596 308956 9648
rect 309008 9636 309014 9648
rect 563238 9636 563244 9648
rect 309008 9608 563244 9636
rect 309008 9596 309014 9608
rect 563238 9596 563244 9608
rect 563296 9596 563302 9648
rect 199930 9528 199936 9580
rect 199988 9568 199994 9580
rect 455690 9568 455696 9580
rect 199988 9540 455696 9568
rect 199988 9528 199994 9540
rect 455690 9528 455696 9540
rect 455748 9528 455754 9580
rect 180242 9460 180248 9512
rect 180300 9500 180306 9512
rect 222838 9500 222844 9512
rect 180300 9472 222844 9500
rect 180300 9460 180306 9472
rect 222838 9460 222844 9472
rect 222896 9460 222902 9512
rect 259270 9460 259276 9512
rect 259328 9500 259334 9512
rect 304350 9500 304356 9512
rect 259328 9472 304356 9500
rect 259328 9460 259334 9472
rect 304350 9460 304356 9472
rect 304408 9460 304414 9512
rect 311802 9460 311808 9512
rect 311860 9500 311866 9512
rect 570322 9500 570328 9512
rect 311860 9472 570328 9500
rect 311860 9460 311866 9472
rect 570322 9460 570328 9472
rect 570380 9460 570386 9512
rect 200022 9392 200028 9444
rect 200080 9432 200086 9444
rect 459186 9432 459192 9444
rect 200080 9404 459192 9432
rect 200080 9392 200086 9404
rect 459186 9392 459192 9404
rect 459244 9392 459250 9444
rect 201402 9324 201408 9376
rect 201460 9364 201466 9376
rect 462774 9364 462780 9376
rect 201460 9336 462780 9364
rect 201460 9324 201466 9336
rect 462774 9324 462780 9336
rect 462832 9324 462838 9376
rect 183738 9256 183744 9308
rect 183796 9296 183802 9308
rect 233326 9296 233332 9308
rect 183796 9268 233332 9296
rect 183796 9256 183802 9268
rect 233326 9256 233332 9268
rect 233384 9256 233390 9308
rect 259362 9256 259368 9308
rect 259420 9296 259426 9308
rect 307938 9296 307944 9308
rect 259420 9268 307944 9296
rect 259420 9256 259426 9268
rect 307938 9256 307944 9268
rect 307996 9256 308002 9308
rect 311710 9256 311716 9308
rect 311768 9296 311774 9308
rect 573910 9296 573916 9308
rect 311768 9268 573916 9296
rect 311768 9256 311774 9268
rect 573910 9256 573916 9268
rect 573968 9256 573974 9308
<<<<<<< HEAD
rect 129642 9188 129648 9240
rect 129700 9228 129706 9240
rect 222194 9228 222200 9240
rect 129700 9200 222200 9228
rect 129700 9188 129706 9200
=======
rect 129550 9188 129556 9240
rect 129608 9228 129614 9240
rect 222194 9228 222200 9240
rect 129608 9200 222200 9228
rect 129608 9188 129614 9200
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 222194 9188 222200 9200
rect 222252 9188 222258 9240
rect 222746 9188 222752 9240
rect 222804 9228 222810 9240
rect 241606 9228 241612 9240
rect 222804 9200 241612 9228
rect 222804 9188 222810 9200
rect 241606 9188 241612 9200
rect 241664 9188 241670 9240
rect 249610 9188 249616 9240
rect 249668 9228 249674 9240
rect 258258 9228 258264 9240
rect 249668 9200 258264 9228
rect 249668 9188 249674 9200
rect 258258 9188 258264 9200
rect 258316 9188 258322 9240
rect 260742 9188 260748 9240
rect 260800 9228 260806 9240
rect 311434 9228 311440 9240
rect 260800 9200 311440 9228
rect 260800 9188 260806 9200
rect 311434 9188 311440 9200
rect 311492 9188 311498 9240
rect 313090 9188 313096 9240
rect 313148 9228 313154 9240
rect 577406 9228 577412 9240
rect 313148 9200 577412 9228
rect 313148 9188 313154 9200
rect 577406 9188 577412 9200
rect 577464 9188 577470 9240
rect 201310 9120 201316 9172
rect 201368 9160 201374 9172
rect 466270 9160 466276 9172
rect 201368 9132 466276 9160
rect 201368 9120 201374 9132
rect 466270 9120 466276 9132
rect 466328 9120 466334 9172
rect 80882 9052 80888 9104
rect 80940 9092 80946 9104
rect 98086 9092 98092 9104
rect 80940 9064 98092 9092
rect 80940 9052 80946 9064
rect 98086 9052 98092 9064
rect 98144 9052 98150 9104
rect 202782 9052 202788 9104
rect 202840 9092 202846 9104
rect 469858 9092 469864 9104
rect 202840 9064 469864 9092
rect 202840 9052 202846 9064
rect 469858 9052 469864 9064
rect 469916 9052 469922 9104
rect 202690 8984 202696 9036
rect 202748 9024 202754 9036
rect 473446 9024 473452 9036
rect 202748 8996 473452 9024
rect 202748 8984 202754 8996
rect 473446 8984 473452 8996
rect 473504 8984 473510 9036
rect 81342 8916 81348 8968
rect 81400 8956 81406 8968
rect 104526 8956 104532 8968
rect 81400 8928 104532 8956
rect 81400 8916 81406 8928
rect 104526 8916 104532 8928
rect 104584 8916 104590 8968
rect 204162 8916 204168 8968
rect 204220 8956 204226 8968
rect 476942 8956 476948 8968
rect 204220 8928 476948 8956
rect 204220 8916 204226 8928
rect 476942 8916 476948 8928
rect 477000 8916 477006 8968
rect 266262 8848 266268 8900
rect 266320 8888 266326 8900
rect 339862 8888 339868 8900
rect 266320 8860 339868 8888
rect 266320 8848 266326 8860
rect 339862 8848 339868 8860
rect 339920 8848 339926 8900
rect 264790 8780 264796 8832
rect 264848 8820 264854 8832
rect 336274 8820 336280 8832
rect 264848 8792 336280 8820
rect 264848 8780 264854 8792
rect 336274 8780 336280 8792
rect 336332 8780 336338 8832
rect 264882 8712 264888 8764
rect 264940 8752 264946 8764
rect 332686 8752 332692 8764
rect 264940 8724 332692 8752
rect 264940 8712 264946 8724
rect 332686 8712 332692 8724
rect 332744 8712 332750 8764
rect 263502 8644 263508 8696
rect 263560 8684 263566 8696
rect 329190 8684 329196 8696
rect 263560 8656 329196 8684
rect 263560 8644 263566 8656
rect 329190 8644 329196 8656
rect 329248 8644 329254 8696
rect 263410 8576 263416 8628
rect 263468 8616 263474 8628
rect 325602 8616 325608 8628
rect 263468 8588 325608 8616
rect 263468 8576 263474 8588
rect 325602 8576 325608 8588
rect 325660 8576 325666 8628
rect 262122 8508 262128 8560
rect 262180 8548 262186 8560
rect 322106 8548 322112 8560
rect 262180 8520 322112 8548
rect 262180 8508 262186 8520
rect 322106 8508 322112 8520
rect 322164 8508 322170 8560
rect 262030 8440 262036 8492
rect 262088 8480 262094 8492
rect 318518 8480 318524 8492
rect 262088 8452 318524 8480
rect 262088 8440 262094 8452
rect 318518 8440 318524 8452
rect 318576 8440 318582 8492
<<<<<<< HEAD
rect 260650 8372 260656 8424
rect 260708 8412 260714 8424
rect 315022 8412 315028 8424
rect 260708 8384 315028 8412
rect 260708 8372 260714 8384
=======
rect 260558 8372 260564 8424
rect 260616 8412 260622 8424
rect 315022 8412 315028 8424
rect 260616 8384 315028 8412
rect 260616 8372 260622 8384
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 315022 8372 315028 8384
rect 315080 8372 315086 8424
rect 184750 8236 184756 8288
rect 184808 8276 184814 8288
rect 384758 8276 384764 8288
rect 184808 8248 384764 8276
rect 184808 8236 184814 8248
rect 384758 8236 384764 8248
rect 384816 8236 384822 8288
rect 186222 8168 186228 8220
rect 186280 8208 186286 8220
rect 388254 8208 388260 8220
rect 186280 8180 388260 8208
rect 186280 8168 186286 8180
rect 388254 8168 388260 8180
rect 388312 8168 388318 8220
rect 187602 8100 187608 8152
rect 187660 8140 187666 8152
rect 391842 8140 391848 8152
rect 187660 8112 391848 8140
rect 187660 8100 187666 8112
rect 391842 8100 391848 8112
rect 391900 8100 391906 8152
rect 187510 8032 187516 8084
rect 187568 8072 187574 8084
rect 395338 8072 395344 8084
rect 187568 8044 395344 8072
rect 187568 8032 187574 8044
rect 395338 8032 395344 8044
rect 395396 8032 395402 8084
rect 188890 7964 188896 8016
rect 188948 8004 188954 8016
rect 398926 8004 398932 8016
rect 188948 7976 398932 8004
rect 188948 7964 188954 7976
rect 398926 7964 398932 7976
rect 398984 7964 398990 8016
rect 188982 7896 188988 7948
rect 189040 7936 189046 7948
rect 402514 7936 402520 7948
rect 189040 7908 402520 7936
rect 189040 7896 189046 7908
rect 402514 7896 402520 7908
rect 402572 7896 402578 7948
rect 190270 7828 190276 7880
rect 190328 7868 190334 7880
rect 406010 7868 406016 7880
rect 190328 7840 406016 7868
rect 190328 7828 190334 7840
rect 406010 7828 406016 7840
rect 406068 7828 406074 7880
rect 411898 7828 411904 7880
rect 411956 7868 411962 7880
rect 480530 7868 480536 7880
rect 411956 7840 480536 7868
rect 411956 7828 411962 7840
rect 480530 7828 480536 7840
rect 480588 7828 480594 7880
rect 190362 7760 190368 7812
rect 190420 7800 190426 7812
rect 409598 7800 409604 7812
rect 190420 7772 409604 7800
rect 190420 7760 190426 7772
rect 409598 7760 409604 7772
rect 409656 7760 409662 7812
rect 410518 7760 410524 7812
rect 410576 7800 410582 7812
rect 495894 7800 495900 7812
rect 410576 7772 495900 7800
rect 410576 7760 410582 7772
rect 495894 7760 495900 7772
rect 495952 7760 495958 7812
rect 191650 7692 191656 7744
rect 191708 7732 191714 7744
rect 413094 7732 413100 7744
rect 191708 7704 413100 7732
rect 191708 7692 191714 7704
rect 413094 7692 413100 7704
rect 413152 7692 413158 7744
rect 413278 7692 413284 7744
rect 413336 7732 413342 7744
rect 505370 7732 505376 7744
rect 413336 7704 505376 7732
rect 413336 7692 413342 7704
rect 505370 7692 505376 7704
rect 505428 7692 505434 7744
rect 83458 7624 83464 7676
rect 83516 7664 83522 7676
rect 93854 7664 93860 7676
rect 83516 7636 93860 7664
rect 83516 7624 83522 7636
rect 93854 7624 93860 7636
rect 93912 7624 93918 7676
rect 191742 7624 191748 7676
rect 191800 7664 191806 7676
rect 416682 7664 416688 7676
rect 191800 7636 416688 7664
rect 191800 7624 191806 7636
rect 416682 7624 416688 7636
rect 416740 7624 416746 7676
rect 418798 7624 418804 7676
rect 418856 7664 418862 7676
rect 492306 7664 492312 7676
rect 418856 7636 492312 7664
rect 418856 7624 418862 7636
rect 492306 7624 492312 7636
rect 492364 7624 492370 7676
rect 51350 7556 51356 7608
rect 51408 7596 51414 7608
rect 69198 7596 69204 7608
rect 51408 7568 69204 7596
rect 51408 7556 51414 7568
rect 69198 7556 69204 7568
rect 69256 7556 69262 7608
rect 70302 7556 70308 7608
rect 70360 7596 70366 7608
rect 94590 7596 94596 7608
rect 70360 7568 94596 7596
rect 70360 7556 70366 7568
rect 94590 7556 94596 7568
rect 94648 7556 94654 7608
rect 106090 7556 106096 7608
rect 106148 7596 106154 7608
rect 116394 7596 116400 7608
rect 106148 7568 116400 7596
rect 106148 7556 106154 7568
rect 116394 7556 116400 7568
rect 116452 7556 116458 7608
rect 193122 7556 193128 7608
rect 193180 7596 193186 7608
rect 420178 7596 420184 7608
rect 193180 7568 420184 7596
rect 193180 7556 193186 7568
rect 420178 7556 420184 7568
rect 420236 7556 420242 7608
rect 184842 7488 184848 7540
rect 184900 7528 184906 7540
rect 381170 7528 381176 7540
rect 184900 7500 381176 7528
rect 184900 7488 184906 7500
rect 381170 7488 381176 7500
rect 381228 7488 381234 7540
rect 183462 7420 183468 7472
rect 183520 7460 183526 7472
rect 377674 7460 377680 7472
rect 183520 7432 377680 7460
rect 183520 7420 183526 7432
rect 377674 7420 377680 7432
rect 377732 7420 377738 7472
rect 183370 7352 183376 7404
rect 183428 7392 183434 7404
rect 374086 7392 374092 7404
rect 183428 7364 374092 7392
rect 183428 7352 183434 7364
rect 374086 7352 374092 7364
rect 374144 7352 374150 7404
rect 181990 7284 181996 7336
rect 182048 7324 182054 7336
rect 370590 7324 370596 7336
rect 182048 7296 370596 7324
rect 182048 7284 182054 7296
rect 370590 7284 370596 7296
rect 370648 7284 370654 7336
rect 371878 7284 371884 7336
rect 371936 7324 371942 7336
rect 487614 7324 487620 7336
rect 371936 7296 487620 7324
rect 371936 7284 371942 7296
rect 487614 7284 487620 7296
rect 487672 7284 487678 7336
rect 182082 7216 182088 7268
rect 182140 7256 182146 7268
rect 367002 7256 367008 7268
rect 182140 7228 367008 7256
rect 182140 7216 182146 7228
rect 367002 7216 367008 7228
rect 367060 7216 367066 7268
rect 180702 7148 180708 7200
rect 180760 7188 180766 7200
rect 363506 7188 363512 7200
rect 180760 7160 363512 7188
rect 180760 7148 180766 7160
rect 363506 7148 363512 7160
rect 363564 7148 363570 7200
rect 180610 7080 180616 7132
rect 180668 7120 180674 7132
rect 359918 7120 359924 7132
rect 180668 7092 359924 7120
rect 180668 7080 180674 7092
rect 359918 7080 359924 7092
rect 359976 7080 359982 7132
rect 179322 7012 179328 7064
rect 179380 7052 179386 7064
rect 356330 7052 356336 7064
rect 179380 7024 356336 7052
rect 179380 7012 179386 7024
rect 356330 7012 356336 7024
rect 356388 7012 356394 7064
rect 206278 6808 206284 6860
rect 206336 6848 206342 6860
rect 232222 6848 232228 6860
rect 206336 6820 232228 6848
rect 206336 6808 206342 6820
rect 232222 6808 232228 6820
rect 232280 6808 232286 6860
rect 255222 6808 255228 6860
rect 255280 6848 255286 6860
rect 283098 6848 283104 6860
rect 255280 6820 283104 6848
rect 255280 6808 255286 6820
rect 283098 6808 283104 6820
rect 283156 6808 283162 6860
rect 302050 6808 302056 6860
rect 302108 6848 302114 6860
rect 527818 6848 527824 6860
rect 302108 6820 527824 6848
rect 302108 6808 302114 6820
rect 527818 6808 527824 6820
rect 527876 6808 527882 6860
rect 205082 6740 205088 6792
rect 205140 6780 205146 6792
rect 237374 6780 237380 6792
rect 205140 6752 237380 6780
rect 205140 6740 205146 6752
rect 237374 6740 237380 6752
rect 237432 6740 237438 6792
rect 255130 6740 255136 6792
rect 255188 6780 255194 6792
rect 286594 6780 286600 6792
rect 255188 6752 286600 6780
rect 255188 6740 255194 6752
rect 286594 6740 286600 6752
rect 286652 6740 286658 6792
rect 303522 6740 303528 6792
rect 303580 6780 303586 6792
rect 531314 6780 531320 6792
rect 303580 6752 531320 6780
rect 303580 6740 303586 6752
rect 531314 6740 531320 6752
rect 531372 6740 531378 6792
rect 204898 6672 204904 6724
rect 204956 6712 204962 6724
rect 239306 6712 239312 6724
rect 204956 6684 239312 6712
rect 204956 6672 204962 6684
rect 239306 6672 239312 6684
rect 239364 6672 239370 6724
rect 256602 6672 256608 6724
rect 256660 6712 256666 6724
rect 290182 6712 290188 6724
rect 256660 6684 290188 6712
rect 256660 6672 256666 6684
rect 290182 6672 290188 6684
rect 290240 6672 290246 6724
rect 303430 6672 303436 6724
rect 303488 6712 303494 6724
rect 534902 6712 534908 6724
rect 303488 6684 534908 6712
rect 303488 6672 303494 6684
rect 534902 6672 534908 6684
rect 534960 6672 534966 6724
rect 155770 6604 155776 6656
rect 155828 6644 155834 6656
rect 235810 6644 235816 6656
rect 155828 6616 235816 6644
rect 155828 6604 155834 6616
rect 235810 6604 235816 6616
rect 235868 6604 235874 6656
rect 237006 6604 237012 6656
rect 237064 6644 237070 6656
rect 244274 6644 244280 6656
rect 237064 6616 244280 6644
rect 237064 6604 237070 6616
rect 244274 6604 244280 6616
rect 244332 6604 244338 6656
rect 256510 6604 256516 6656
rect 256568 6644 256574 6656
rect 293678 6644 293684 6656
rect 256568 6616 293684 6644
rect 256568 6604 256574 6616
rect 293678 6604 293684 6616
rect 293736 6604 293742 6656
rect 304810 6604 304816 6656
rect 304868 6644 304874 6656
rect 538398 6644 538404 6656
rect 304868 6616 538404 6644
rect 304868 6604 304874 6616
rect 538398 6604 538404 6616
rect 538456 6604 538462 6656
rect 157242 6536 157248 6588
rect 157300 6576 157306 6588
rect 242894 6576 242900 6588
rect 157300 6548 242900 6576
rect 157300 6536 157306 6548
rect 242894 6536 242900 6548
rect 242952 6536 242958 6588
rect 257890 6536 257896 6588
rect 257948 6576 257954 6588
rect 297266 6576 297272 6588
rect 257948 6548 297272 6576
rect 257948 6536 257954 6548
rect 297266 6536 297272 6548
rect 297324 6536 297330 6588
rect 304902 6536 304908 6588
rect 304960 6576 304966 6588
rect 541986 6576 541992 6588
rect 304960 6548 541992 6576
rect 304960 6536 304966 6548
rect 541986 6536 541992 6548
rect 542044 6536 542050 6588
rect 79318 6468 79324 6520
rect 79376 6508 79382 6520
rect 90358 6508 90364 6520
rect 79376 6480 90364 6508
rect 79376 6468 79382 6480
rect 90358 6468 90364 6480
rect 90416 6468 90422 6520
rect 160002 6468 160008 6520
rect 160060 6508 160066 6520
rect 257062 6508 257068 6520
rect 160060 6480 257068 6508
rect 160060 6468 160066 6480
rect 257062 6468 257068 6480
rect 257120 6468 257126 6520
rect 257982 6468 257988 6520
rect 258040 6508 258046 6520
rect 300762 6508 300768 6520
rect 258040 6480 300768 6508
rect 258040 6468 258046 6480
rect 300762 6468 300768 6480
rect 300820 6468 300826 6520
rect 306190 6468 306196 6520
rect 306248 6508 306254 6520
rect 545482 6508 545488 6520
rect 306248 6480 545488 6508
rect 306248 6468 306254 6480
rect 545482 6468 545488 6480
rect 545540 6468 545546 6520
rect 167178 6400 167184 6452
rect 167236 6440 167242 6452
rect 289078 6440 289084 6452
rect 167236 6412 289084 6440
rect 167236 6400 167242 6412
rect 289078 6400 289084 6412
rect 289136 6400 289142 6452
rect 306282 6400 306288 6452
rect 306340 6440 306346 6452
rect 549070 6440 549076 6452
rect 306340 6412 549076 6440
rect 306340 6400 306346 6412
rect 549070 6400 549076 6412
rect 549128 6400 549134 6452
rect 42794 6332 42800 6384
rect 42852 6372 42858 6384
rect 89898 6372 89904 6384
rect 42852 6344 89904 6372
rect 42852 6332 42858 6344
rect 89898 6332 89904 6344
rect 89956 6332 89962 6384
rect 166810 6332 166816 6384
rect 166868 6372 166874 6384
rect 288986 6372 288992 6384
rect 166868 6344 288992 6372
rect 166868 6332 166874 6344
rect 288986 6332 288992 6344
rect 289044 6332 289050 6384
rect 307662 6332 307668 6384
rect 307720 6372 307726 6384
rect 552658 6372 552664 6384
rect 307720 6344 552664 6372
rect 307720 6332 307726 6344
rect 552658 6332 552664 6344
rect 552716 6332 552722 6384
rect 34790 6264 34796 6316
rect 34848 6304 34854 6316
rect 88334 6304 88340 6316
rect 34848 6276 88340 6304
rect 34848 6264 34854 6276
rect 88334 6264 88340 6276
rect 88392 6264 88398 6316
rect 166902 6264 166908 6316
rect 166960 6304 166966 6316
rect 292574 6304 292580 6316
rect 166960 6276 292580 6304
rect 166960 6264 166966 6276
rect 292574 6264 292580 6276
rect 292632 6264 292638 6316
rect 307570 6264 307576 6316
rect 307628 6304 307634 6316
rect 556154 6304 556160 6316
rect 307628 6276 556160 6304
rect 307628 6264 307634 6276
rect 556154 6264 556160 6276
rect 556212 6264 556218 6316
rect 2866 6196 2872 6248
rect 2924 6236 2930 6248
rect 57238 6236 57244 6248
rect 2924 6208 57244 6236
rect 2924 6196 2930 6208
rect 57238 6196 57244 6208
rect 57296 6196 57302 6248
rect 63218 6196 63224 6248
rect 63276 6236 63282 6248
rect 93946 6236 93952 6248
rect 63276 6208 93952 6236
rect 63276 6196 63282 6208
rect 93946 6196 93952 6208
rect 94004 6196 94010 6248
rect 168282 6196 168288 6248
rect 168340 6236 168346 6248
rect 296070 6236 296076 6248
rect 168340 6208 296076 6236
rect 168340 6196 168346 6208
rect 296070 6196 296076 6208
rect 296128 6196 296134 6248
rect 309042 6196 309048 6248
rect 309100 6236 309106 6248
rect 559742 6236 559748 6248
rect 309100 6208 559748 6236
rect 309100 6196 309106 6208
rect 559742 6196 559748 6208
rect 559800 6196 559806 6248
rect 27706 6128 27712 6180
rect 27764 6168 27770 6180
rect 86954 6168 86960 6180
rect 27764 6140 86960 6168
rect 27764 6128 27770 6140
rect 86954 6128 86960 6140
rect 87012 6128 87018 6180
rect 87966 6128 87972 6180
rect 88024 6168 88030 6180
rect 98638 6168 98644 6180
rect 88024 6140 98644 6168
rect 88024 6128 88030 6140
rect 98638 6128 98644 6140
rect 98696 6128 98702 6180
rect 141878 6128 141884 6180
rect 141936 6168 141942 6180
rect 164878 6168 164884 6180
rect 141936 6140 164884 6168
rect 141936 6128 141942 6140
rect 164878 6128 164884 6140
rect 164936 6128 164942 6180
rect 168190 6128 168196 6180
rect 168248 6168 168254 6180
rect 299658 6168 299664 6180
rect 168248 6140 299664 6168
rect 168248 6128 168254 6140
rect 299658 6128 299664 6140
rect 299716 6128 299722 6180
rect 310422 6128 310428 6180
rect 310480 6168 310486 6180
rect 566826 6168 566832 6180
rect 310480 6140 566832 6168
rect 310480 6128 310486 6140
rect 566826 6128 566832 6140
rect 566884 6128 566890 6180
rect 204990 6060 204996 6112
rect 205048 6100 205054 6112
rect 228726 6100 228732 6112
rect 205048 6072 228732 6100
rect 205048 6060 205054 6072
rect 228726 6060 228732 6072
rect 228784 6060 228790 6112
rect 229830 6060 229836 6112
rect 229888 6100 229894 6112
rect 242158 6100 242164 6112
rect 229888 6072 242164 6100
rect 229888 6060 229894 6072
rect 242158 6060 242164 6072
rect 242216 6060 242222 6112
rect 253750 6060 253756 6112
rect 253808 6100 253814 6112
rect 279510 6100 279516 6112
rect 253808 6072 279516 6100
rect 253808 6060 253814 6072
rect 279510 6060 279516 6072
rect 279568 6060 279574 6112
rect 302142 6060 302148 6112
rect 302200 6100 302206 6112
rect 524230 6100 524236 6112
rect 302200 6072 524236 6100
rect 302200 6060 302206 6072
rect 524230 6060 524236 6072
rect 524288 6060 524294 6112
rect 224218 5992 224224 6044
rect 224276 6032 224282 6044
rect 246390 6032 246396 6044
rect 224276 6004 246396 6032
rect 224276 5992 224282 6004
rect 246390 5992 246396 6004
rect 246448 5992 246454 6044
rect 253842 5992 253848 6044
rect 253900 6032 253906 6044
rect 276014 6032 276020 6044
rect 253900 6004 276020 6032
rect 253900 5992 253906 6004
rect 276014 5992 276020 6004
rect 276072 5992 276078 6044
rect 300670 5992 300676 6044
rect 300728 6032 300734 6044
rect 520734 6032 520740 6044
rect 300728 6004 520740 6032
rect 300728 5992 300734 6004
rect 520734 5992 520740 6004
rect 520792 5992 520798 6044
rect 219250 5924 219256 5976
rect 219308 5964 219314 5976
rect 240134 5964 240140 5976
rect 219308 5936 240140 5964
rect 219308 5924 219314 5936
rect 240134 5924 240140 5936
rect 240192 5924 240198 5976
rect 252370 5924 252376 5976
rect 252428 5964 252434 5976
rect 272426 5964 272432 5976
rect 252428 5936 272432 5964
rect 252428 5924 252434 5936
rect 272426 5924 272432 5936
rect 272484 5924 272490 5976
rect 300578 5924 300584 5976
rect 300636 5964 300642 5976
rect 517146 5964 517152 5976
rect 300636 5936 517152 5964
rect 300636 5924 300642 5936
rect 517146 5924 517152 5936
rect 517204 5924 517210 5976
rect 212166 5856 212172 5908
rect 212224 5896 212230 5908
rect 231118 5896 231124 5908
rect 212224 5868 231124 5896
rect 212224 5856 212230 5868
rect 231118 5856 231124 5868
rect 231176 5856 231182 5908
rect 251082 5856 251088 5908
rect 251140 5896 251146 5908
rect 261754 5896 261760 5908
rect 251140 5868 261760 5896
rect 251140 5856 251146 5868
rect 261754 5856 261760 5868
rect 261812 5856 261818 5908
rect 299198 5856 299204 5908
rect 299256 5896 299262 5908
rect 513558 5896 513564 5908
rect 299256 5868 513564 5896
rect 299256 5856 299262 5868
rect 513558 5856 513564 5868
rect 513616 5856 513622 5908
rect 299290 5788 299296 5840
rect 299348 5828 299354 5840
rect 510062 5828 510068 5840
rect 299348 5800 510068 5828
rect 299348 5788 299354 5800
rect 510062 5788 510068 5800
rect 510120 5788 510126 5840
rect 297910 5720 297916 5772
rect 297968 5760 297974 5772
<<<<<<< HEAD
rect 506566 5760 506572 5772
rect 297968 5732 506572 5760
rect 297968 5720 297974 5732
rect 506566 5720 506572 5732
rect 506624 5720 506630 5772
=======
rect 506474 5760 506480 5772
rect 297968 5732 506480 5760
rect 297968 5720 297974 5732
rect 506474 5720 506480 5732
rect 506532 5720 506538 5772
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 298002 5652 298008 5704
rect 298060 5692 298066 5704
rect 502978 5692 502984 5704
rect 298060 5664 502984 5692
rect 298060 5652 298066 5664
rect 502978 5652 502984 5664
rect 503036 5652 503042 5704
rect 406378 5584 406384 5636
rect 406436 5624 406442 5636
rect 580166 5624 580172 5636
rect 406436 5596 580172 5624
rect 406436 5584 406442 5596
rect 580166 5584 580172 5596
rect 580224 5584 580230 5636
rect 69106 5516 69112 5568
rect 69164 5556 69170 5568
rect 72418 5556 72424 5568
rect 69164 5528 72424 5556
rect 69164 5516 69170 5528
rect 72418 5516 72424 5528
rect 72476 5516 72482 5568
rect 98638 5516 98644 5568
rect 98696 5556 98702 5568
rect 100754 5556 100760 5568
rect 98696 5528 100760 5556
rect 98696 5516 98702 5528
rect 100754 5516 100760 5528
rect 100812 5516 100818 5568
rect 104710 5516 104716 5568
rect 104768 5556 104774 5568
rect 112806 5556 112812 5568
rect 104768 5528 112812 5556
rect 104768 5516 104774 5528
rect 112806 5516 112812 5528
rect 112864 5516 112870 5568
rect 244090 5516 244096 5568
rect 244148 5556 244154 5568
rect 245654 5556 245660 5568
rect 244148 5528 245660 5556
rect 244148 5516 244154 5528
rect 245654 5516 245660 5528
rect 245712 5516 245718 5568
rect 246942 5516 246948 5568
rect 247000 5556 247006 5568
rect 247586 5556 247592 5568
rect 247000 5528 247592 5556
rect 247000 5516 247006 5528
rect 247586 5516 247592 5528
rect 247644 5516 247650 5568
rect 249702 5516 249708 5568
rect 249760 5556 249766 5568
rect 254670 5556 254676 5568
rect 249760 5528 254676 5556
rect 249760 5516 249766 5528
rect 254670 5516 254676 5528
rect 254728 5516 254734 5568
rect 146202 5448 146208 5500
rect 146260 5488 146266 5500
rect 186130 5488 186136 5500
rect 146260 5460 186136 5488
rect 146260 5448 146266 5460
rect 186130 5448 186136 5460
rect 186188 5448 186194 5500
rect 215202 5448 215208 5500
rect 215260 5488 215266 5500
rect 537202 5488 537208 5500
rect 215260 5460 537208 5488
rect 215260 5448 215266 5460
rect 537202 5448 537208 5460
rect 537260 5448 537266 5500
rect 79962 5380 79968 5432
rect 80020 5420 80026 5432
rect 97442 5420 97448 5432
rect 80020 5392 97448 5420
rect 80020 5380 80026 5392
rect 97442 5380 97448 5392
rect 97500 5380 97506 5432
rect 147582 5380 147588 5432
rect 147640 5420 147646 5432
rect 189718 5420 189724 5432
rect 147640 5392 189724 5420
rect 147640 5380 147646 5392
rect 189718 5380 189724 5392
rect 189776 5380 189782 5432
rect 216490 5380 216496 5432
rect 216548 5420 216554 5432
rect 540790 5420 540796 5432
rect 216548 5392 540796 5420
rect 216548 5380 216554 5392
rect 540790 5380 540796 5392
rect 540848 5380 540854 5432
rect 84470 5312 84476 5364
rect 84528 5352 84534 5364
rect 97994 5352 98000 5364
rect 84528 5324 98000 5352
rect 84528 5312 84534 5324
rect 97994 5312 98000 5324
rect 98052 5312 98058 5364
rect 147490 5312 147496 5364
rect 147548 5352 147554 5364
rect 193214 5352 193220 5364
rect 147548 5324 193220 5352
rect 147548 5312 147554 5324
rect 193214 5312 193220 5324
rect 193272 5312 193278 5364
rect 216582 5312 216588 5364
rect 216640 5352 216646 5364
rect 544378 5352 544384 5364
rect 216640 5324 544384 5352
rect 216640 5312 216646 5324
rect 544378 5312 544384 5324
rect 544436 5312 544442 5364
rect 77386 5244 77392 5296
rect 77444 5284 77450 5296
rect 96798 5284 96804 5296
rect 77444 5256 96804 5284
rect 77444 5244 77450 5256
rect 96798 5244 96804 5256
rect 96856 5244 96862 5296
rect 148870 5244 148876 5296
rect 148928 5284 148934 5296
rect 196802 5284 196808 5296
rect 148928 5256 196808 5284
rect 148928 5244 148934 5256
rect 196802 5244 196808 5256
rect 196860 5244 196866 5296
rect 217870 5244 217876 5296
rect 217928 5284 217934 5296
rect 547874 5284 547880 5296
rect 217928 5256 547880 5284
rect 217928 5244 217934 5256
rect 547874 5244 547880 5256
rect 547932 5244 547938 5296
rect 79870 5176 79876 5228
rect 79928 5216 79934 5228
rect 101030 5216 101036 5228
rect 79928 5188 101036 5216
rect 79928 5176 79934 5188
rect 101030 5176 101036 5188
rect 101088 5176 101094 5228
rect 148778 5176 148784 5228
rect 148836 5216 148842 5228
rect 200298 5216 200304 5228
rect 148836 5188 200304 5216
rect 148836 5176 148842 5188
rect 200298 5176 200304 5188
rect 200356 5176 200362 5228
rect 217962 5176 217968 5228
rect 218020 5216 218026 5228
rect 551462 5216 551468 5228
rect 218020 5188 551468 5216
rect 218020 5176 218026 5188
rect 551462 5176 551468 5188
rect 551520 5176 551526 5228
rect 52546 5108 52552 5160
rect 52604 5148 52610 5160
rect 65518 5148 65524 5160
rect 52604 5120 65524 5148
rect 52604 5108 52610 5120
rect 65518 5108 65524 5120
rect 65576 5108 65582 5160
rect 73798 5108 73804 5160
rect 73856 5148 73862 5160
rect 96706 5148 96712 5160
rect 73856 5120 96712 5148
rect 73856 5108 73862 5120
rect 96706 5108 96712 5120
rect 96764 5108 96770 5160
rect 150250 5108 150256 5160
rect 150308 5148 150314 5160
rect 203886 5148 203892 5160
rect 150308 5120 203892 5148
rect 150308 5108 150314 5120
rect 203886 5108 203892 5120
rect 203944 5108 203950 5160
rect 219158 5108 219164 5160
rect 219216 5148 219222 5160
rect 554958 5148 554964 5160
rect 219216 5120 554964 5148
rect 219216 5108 219222 5120
rect 554958 5108 554964 5120
rect 555016 5108 555022 5160
rect 44266 5040 44272 5092
rect 44324 5080 44330 5092
rect 67726 5080 67732 5092
rect 44324 5052 67732 5080
rect 44324 5040 44330 5052
rect 67726 5040 67732 5052
rect 67784 5040 67790 5092
rect 77202 5040 77208 5092
rect 77260 5080 77266 5092
rect 85758 5080 85764 5092
rect 77260 5052 85764 5080
rect 77260 5040 77266 5052
rect 85758 5040 85764 5052
rect 85816 5040 85822 5092
rect 86218 5040 86224 5092
rect 86276 5080 86282 5092
rect 111610 5080 111616 5092
rect 86276 5052 111616 5080
rect 86276 5040 86282 5052
rect 111610 5040 111616 5052
rect 111668 5040 111674 5092
rect 150342 5040 150348 5092
rect 150400 5080 150406 5092
rect 207382 5080 207388 5092
rect 150400 5052 207388 5080
rect 150400 5040 150406 5052
rect 207382 5040 207388 5052
rect 207440 5040 207446 5092
rect 219342 5040 219348 5092
rect 219400 5080 219406 5092
rect 558546 5080 558552 5092
rect 219400 5052 558552 5080
rect 219400 5040 219406 5052
rect 558546 5040 558552 5052
rect 558604 5040 558610 5092
rect 21818 4972 21824 5024
rect 21876 5012 21882 5024
rect 53098 5012 53104 5024
rect 21876 4984 53104 5012
rect 21876 4972 21882 4984
rect 53098 4972 53104 4984
rect 53156 4972 53162 5024
rect 59630 4972 59636 5024
rect 59688 5012 59694 5024
rect 93118 5012 93124 5024
rect 59688 4984 93124 5012
rect 59688 4972 59694 4984
rect 93118 4972 93124 4984
rect 93176 4972 93182 5024
rect 151722 4972 151728 5024
rect 151780 5012 151786 5024
rect 210970 5012 210976 5024
rect 151780 4984 210976 5012
rect 151780 4972 151786 4984
rect 210970 4972 210976 4984
rect 211028 4972 211034 5024
rect 220630 4972 220636 5024
rect 220688 5012 220694 5024
rect 562042 5012 562048 5024
rect 220688 4984 562048 5012
rect 220688 4972 220694 4984
rect 562042 4972 562048 4984
rect 562100 4972 562106 5024
rect 4062 4904 4068 4956
rect 4120 4944 4126 4956
rect 50338 4944 50344 4956
rect 4120 4916 50344 4944
rect 4120 4904 4126 4916
rect 50338 4904 50344 4916
rect 50396 4904 50402 4956
rect 56042 4904 56048 4956
rect 56100 4944 56106 4956
rect 92566 4944 92572 4956
rect 56100 4916 92572 4944
rect 56100 4904 56106 4916
rect 92566 4904 92572 4916
rect 92624 4904 92630 4956
rect 106182 4904 106188 4956
rect 106240 4944 106246 4956
rect 116486 4944 116492 4956
rect 106240 4916 116492 4944
rect 106240 4904 106246 4916
rect 116486 4904 116492 4916
rect 116544 4904 116550 4956
rect 151630 4904 151636 4956
rect 151688 4944 151694 4956
rect 214466 4944 214472 4956
rect 151688 4916 214472 4944
rect 151688 4904 151694 4916
rect 214466 4904 214472 4916
rect 214524 4904 214530 4956
rect 220722 4904 220728 4956
rect 220780 4944 220786 4956
rect 565630 4944 565636 4956
rect 220780 4916 565636 4944
rect 220780 4904 220786 4916
rect 565630 4904 565636 4916
rect 565688 4904 565694 4956
rect 7650 4836 7656 4888
rect 7708 4876 7714 4888
rect 60826 4876 60832 4888
rect 7708 4848 60832 4876
rect 7708 4836 7714 4848
rect 60826 4836 60832 4848
rect 60884 4836 60890 4888
rect 62022 4836 62028 4888
rect 62080 4876 62086 4888
rect 69658 4876 69664 4888
rect 62080 4848 69664 4876
rect 62080 4836 62086 4848
rect 69658 4836 69664 4848
rect 69716 4836 69722 4888
rect 84102 4836 84108 4888
rect 84160 4876 84166 4888
rect 118786 4876 118792 4888
rect 84160 4848 118792 4876
rect 84160 4836 84166 4848
rect 118786 4836 118792 4848
rect 118844 4836 118850 4888
rect 153010 4836 153016 4888
rect 153068 4876 153074 4888
rect 218054 4876 218060 4888
rect 153068 4848 218060 4876
rect 153068 4836 153074 4848
rect 218054 4836 218060 4848
rect 218112 4836 218118 4888
rect 222102 4836 222108 4888
rect 222160 4876 222166 4888
rect 569126 4876 569132 4888
rect 222160 4848 569132 4876
rect 222160 4836 222166 4848
rect 569126 4836 569132 4848
rect 569184 4836 569190 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 58618 4808 58624 4820
rect 624 4780 58624 4808
rect 624 4768 630 4780
rect 58618 4768 58624 4780
rect 58676 4768 58682 4820
rect 84010 4768 84016 4820
rect 84068 4808 84074 4820
rect 122282 4808 122288 4820
rect 84068 4780 122288 4808
rect 84068 4768 84074 4780
rect 122282 4768 122288 4780
rect 122340 4768 122346 4820
rect 153102 4768 153108 4820
rect 153160 4808 153166 4820
rect 221550 4808 221556 4820
rect 153160 4780 221556 4808
rect 153160 4768 153166 4780
rect 221550 4768 221556 4780
rect 221608 4768 221614 4820
rect 222010 4768 222016 4820
rect 222068 4808 222074 4820
rect 572714 4808 572720 4820
rect 222068 4780 572720 4808
rect 222068 4768 222074 4780
rect 572714 4768 572720 4780
rect 572772 4768 572778 4820
rect 58434 4700 58440 4752
rect 58492 4740 58498 4752
rect 70578 4740 70584 4752
rect 58492 4712 70584 4740
rect 58492 4700 58498 4712
rect 70578 4700 70584 4712
rect 70636 4700 70642 4752
rect 146110 4700 146116 4752
rect 146168 4740 146174 4752
rect 182542 4740 182548 4752
rect 146168 4712 182548 4740
rect 146168 4700 146174 4712
rect 182542 4700 182548 4712
rect 182600 4700 182606 4752
rect 215110 4700 215116 4752
rect 215168 4740 215174 4752
rect 533706 4740 533712 4752
rect 215168 4712 533712 4740
rect 215168 4700 215174 4712
rect 533706 4700 533712 4712
rect 533764 4700 533770 4752
rect 144638 4632 144644 4684
rect 144696 4672 144702 4684
rect 179046 4672 179052 4684
rect 144696 4644 179052 4672
rect 144696 4632 144702 4644
rect 179046 4632 179052 4644
rect 179104 4632 179110 4684
rect 213730 4632 213736 4684
rect 213788 4672 213794 4684
rect 530118 4672 530124 4684
rect 213788 4644 530124 4672
rect 213788 4632 213794 4644
rect 530118 4632 530124 4644
rect 530176 4632 530182 4684
rect 144546 4564 144552 4616
rect 144604 4604 144610 4616
rect 175458 4604 175464 4616
rect 144604 4576 175464 4604
rect 144604 4564 144610 4576
rect 175458 4564 175464 4576
rect 175516 4564 175522 4616
rect 213822 4564 213828 4616
rect 213880 4604 213886 4616
rect 526622 4604 526628 4616
rect 213880 4576 526628 4604
rect 213880 4564 213886 4576
rect 526622 4564 526628 4576
rect 526680 4564 526686 4616
rect 91554 4496 91560 4548
rect 91612 4536 91618 4548
rect 94498 4536 94504 4548
rect 91612 4508 94504 4536
rect 91612 4496 91618 4508
rect 94498 4496 94504 4508
rect 94556 4496 94562 4548
rect 143350 4496 143356 4548
rect 143408 4536 143414 4548
rect 171962 4536 171968 4548
rect 143408 4508 171968 4536
rect 143408 4496 143414 4508
rect 171962 4496 171968 4508
rect 172020 4496 172026 4548
rect 212442 4496 212448 4548
rect 212500 4536 212506 4548
rect 523034 4536 523040 4548
rect 212500 4508 523040 4536
rect 212500 4496 212506 4508
rect 523034 4496 523040 4508
rect 523092 4496 523098 4548
rect 143442 4428 143448 4480
rect 143500 4468 143506 4480
rect 168374 4468 168380 4480
rect 143500 4440 168380 4468
rect 143500 4428 143506 4440
rect 168374 4428 168380 4440
rect 168432 4428 168438 4480
rect 212350 4428 212356 4480
rect 212408 4468 212414 4480
rect 519538 4468 519544 4480
rect 212408 4440 519544 4468
rect 212408 4428 212414 4440
rect 519538 4428 519544 4440
rect 519596 4428 519602 4480
rect 211062 4360 211068 4412
rect 211120 4400 211126 4412
rect 515950 4400 515956 4412
rect 211120 4372 515956 4400
rect 211120 4360 211126 4372
rect 515950 4360 515956 4372
rect 516008 4360 516014 4412
rect 210878 4292 210884 4344
rect 210936 4332 210942 4344
rect 512454 4332 512460 4344
rect 210936 4304 512460 4332
rect 210936 4292 210942 4304
rect 512454 4292 512460 4304
rect 512512 4292 512518 4344
rect 65518 4224 65524 4276
rect 65576 4264 65582 4276
rect 71958 4264 71964 4276
rect 65576 4236 71964 4264
rect 65576 4224 65582 4236
rect 71958 4224 71964 4236
rect 72016 4224 72022 4276
rect 75822 4224 75828 4276
rect 75880 4264 75886 4276
rect 79686 4264 79692 4276
rect 75880 4236 79692 4264
rect 75880 4224 75886 4236
rect 79686 4224 79692 4236
rect 79744 4224 79750 4276
<<<<<<< HEAD
rect 103793 4267 103851 4273
rect 103793 4233 103805 4267
rect 103839 4264 103851 4267
rect 109218 4264 109224 4276
rect 103839 4236 109224 4264
rect 103839 4233 103851 4236
rect 103793 4227 103851 4233
rect 109218 4224 109224 4236
rect 109276 4224 109282 4276
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 154482 4224 154488 4276
rect 154540 4264 154546 4276
rect 225138 4264 225144 4276
rect 154540 4236 225144 4264
rect 154540 4224 154546 4236
rect 225138 4224 225144 4236
rect 225196 4224 225202 4276
<<<<<<< HEAD
rect 268838 4264 268844 4276
rect 258046 4236 268844 4264
=======
rect 252462 4224 252468 4276
rect 252520 4264 252526 4276
rect 268838 4264 268844 4276
rect 252520 4236 268844 4264
rect 252520 4224 252526 4236
rect 268838 4224 268844 4236
rect 268896 4224 268902 4276
rect 269022 4224 269028 4276
rect 269080 4264 269086 4276
rect 354030 4264 354036 4276
rect 269080 4236 354036 4264
rect 269080 4224 269086 4236
rect 354030 4224 354036 4236
rect 354088 4224 354094 4276
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 48958 4156 48964 4208
rect 49016 4196 49022 4208
rect 51718 4196 51724 4208
rect 49016 4168 51724 4196
rect 49016 4156 49022 4168
rect 51718 4156 51724 4168
rect 51776 4156 51782 4208
rect 66714 4156 66720 4208
rect 66772 4196 66778 4208
rect 68278 4196 68284 4208
rect 66772 4168 68284 4196
rect 66772 4156 66778 4168
rect 68278 4156 68284 4168
rect 68336 4156 68342 4208
rect 75730 4156 75736 4208
rect 75788 4196 75794 4208
rect 76190 4196 76196 4208
rect 75788 4168 76196 4196
rect 75788 4156 75794 4168
rect 76190 4156 76196 4168
rect 76248 4156 76254 4208
rect 77110 4156 77116 4208
rect 77168 4196 77174 4208
rect 83274 4196 83280 4208
rect 77168 4168 83280 4196
rect 77168 4156 77174 4168
rect 83274 4156 83280 4168
rect 83332 4156 83338 4208
rect 85758 4156 85764 4208
rect 85816 4196 85822 4208
rect 86862 4196 86868 4208
rect 85816 4168 86868 4196
rect 85816 4156 85822 4168
rect 86862 4156 86868 4168
rect 86920 4156 86926 4208
rect 95142 4156 95148 4208
rect 95200 4196 95206 4208
rect 100938 4196 100944 4208
rect 95200 4168 100944 4196
rect 95200 4156 95206 4168
rect 100938 4156 100944 4168
rect 100996 4156 101002 4208
rect 104802 4156 104808 4208
rect 104860 4196 104866 4208
rect 109310 4196 109316 4208
rect 104860 4168 109316 4196
rect 104860 4156 104866 4168
rect 109310 4156 109316 4168
rect 109368 4156 109374 4208
rect 194410 4156 194416 4208
rect 194468 4196 194474 4208
rect 197998 4196 198004 4208
rect 194468 4168 198004 4196
rect 194468 4156 194474 4168
rect 197998 4156 198004 4168
rect 198056 4156 198062 4208
<<<<<<< HEAD
rect 252462 4156 252468 4208
rect 252520 4196 252526 4208
rect 258046 4196 258074 4236
rect 268838 4224 268844 4236
rect 268896 4224 268902 4276
rect 269022 4224 269028 4276
rect 269080 4264 269086 4276
rect 354030 4264 354036 4276
rect 269080 4236 354036 4264
rect 269080 4224 269086 4236
rect 354030 4224 354036 4236
rect 354088 4224 354094 4276
rect 252520 4168 258074 4196
rect 252520 4156 252526 4168
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 472618 4156 472624 4208
rect 472676 4196 472682 4208
rect 474550 4196 474556 4208
rect 472676 4168 474556 4196
rect 472676 4156 472682 4168
rect 474550 4156 474556 4168
rect 474608 4156 474614 4208
rect 64322 4088 64328 4140
rect 64380 4128 64386 4140
rect 116026 4128 116032 4140
rect 64380 4100 116032 4128
rect 64380 4088 64386 4100
rect 116026 4088 116032 4100
rect 116084 4088 116090 4140
<<<<<<< HEAD
rect 137738 4088 137744 4140
rect 137796 4128 137802 4140
rect 143534 4128 143540 4140
rect 137796 4100 143540 4128
rect 137796 4088 137802 4100
rect 143534 4088 143540 4100
rect 143592 4088 143598 4140
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 266538 4088 266544 4140
rect 266596 4128 266602 4140
rect 339586 4128 339592 4140
rect 266596 4100 339592 4128
rect 266596 4088 266602 4100
rect 339586 4088 339592 4100
rect 339644 4088 339650 4140
rect 361390 4088 361396 4140
rect 361448 4128 361454 4140
rect 372890 4128 372896 4140
rect 361448 4100 372896 4128
rect 361448 4088 361454 4100
rect 372890 4088 372896 4100
rect 372948 4088 372954 4140
rect 379422 4088 379428 4140
rect 379480 4128 379486 4140
rect 465166 4128 465172 4140
rect 379480 4100 465172 4128
rect 379480 4088 379486 4100
rect 465166 4088 465172 4100
rect 465224 4088 465230 4140
rect 60826 4020 60832 4072
rect 60884 4060 60890 4072
rect 116118 4060 116124 4072
rect 60884 4032 116124 4060
rect 60884 4020 60890 4032
rect 116118 4020 116124 4032
rect 116176 4020 116182 4072
rect 216858 4020 216864 4072
rect 216916 4060 216922 4072
rect 227070 4060 227076 4072
rect 216916 4032 227076 4060
rect 216916 4020 216922 4032
rect 227070 4020 227076 4032
rect 227128 4020 227134 4072
rect 262950 4020 262956 4072
rect 263008 4060 263014 4072
rect 338114 4060 338120 4072
rect 263008 4032 338120 4060
rect 263008 4020 263014 4032
rect 338114 4020 338120 4032
rect 338172 4020 338178 4072
<<<<<<< HEAD
rect 344554 4020 344560 4072
rect 344612 4060 344618 4072
rect 354674 4060 354680 4072
rect 344612 4032 354680 4060
rect 344612 4020 344618 4032
rect 354674 4020 354680 4032
rect 354732 4020 354738 4072
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 380802 4020 380808 4072
rect 380860 4060 380866 4072
rect 472250 4060 472256 4072
rect 380860 4032 472256 4060
rect 380860 4020 380866 4032
rect 472250 4020 472256 4032
rect 472308 4020 472314 4072
rect 14734 3952 14740 4004
rect 14792 3992 14798 4004
rect 18598 3992 18604 4004
rect 14792 3964 18604 3992
rect 14792 3952 14798 3964
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 57238 3952 57244 4004
rect 57296 3992 57302 4004
<<<<<<< HEAD
rect 103977 3995 104035 4001
rect 103977 3992 103989 3995
rect 57296 3964 103989 3992
rect 57296 3952 57302 3964
rect 103977 3961 103989 3964
rect 104023 3961 104035 3995
rect 103977 3955 104035 3961
rect 105633 3995 105691 4001
rect 105633 3961 105645 3995
rect 105679 3992 105691 3995
rect 107746 3992 107752 4004
rect 105679 3964 107752 3992
rect 105679 3961 105691 3964
rect 105633 3955 105691 3961
rect 107746 3952 107752 3964
rect 107804 3952 107810 4004
=======
rect 108301 3995 108359 4001
rect 108301 3992 108313 3995
rect 57296 3964 108313 3992
rect 57296 3952 57302 3964
rect 108301 3961 108313 3964
rect 108347 3961 108359 3995
rect 108301 3955 108359 3961
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 188522 3952 188528 4004
rect 188580 3992 188586 4004
rect 195238 3992 195244 4004
rect 188580 3964 195244 3992
rect 188580 3952 188586 3964
rect 195238 3952 195244 3964
rect 195296 3952 195302 4004
rect 223942 3952 223948 4004
rect 224000 3992 224006 4004
rect 238018 3992 238024 4004
rect 224000 3964 238024 3992
rect 224000 3952 224006 3964
rect 238018 3952 238024 3964
rect 238076 3952 238082 4004
<<<<<<< HEAD
rect 259546 3952 259552 4004
rect 259604 3992 259610 4004
rect 338390 3992 338396 4004
rect 259604 3964 338396 3992
rect 259604 3952 259610 3964
rect 338390 3952 338396 3964
rect 338448 3952 338454 4004
rect 352006 3992 352012 4004
rect 345676 3964 352012 3992
=======
rect 259454 3952 259460 4004
rect 259512 3992 259518 4004
rect 338390 3992 338396 4004
rect 259512 3964 338396 3992
rect 259512 3952 259518 3964
rect 338390 3952 338396 3964
rect 338448 3952 338454 4004
rect 344554 3952 344560 4004
rect 344612 3992 344618 4004
rect 354674 3992 354680 4004
rect 344612 3964 354680 3992
rect 344612 3952 344618 3964
rect 354674 3952 354680 3964
rect 354732 3952 354738 4004
rect 361482 3952 361488 4004
rect 361540 3992 361546 4004
rect 376478 3992 376484 4004
rect 361540 3964 376484 3992
rect 361540 3952 361546 3964
rect 376478 3952 376484 3964
rect 376536 3952 376542 4004
rect 382182 3952 382188 4004
rect 382240 3992 382246 4004
rect 479334 3992 479340 4004
rect 382240 3964 479340 3992
rect 382240 3952 382246 3964
rect 479334 3952 479340 3964
rect 479392 3952 479398 4004
rect 489914 3952 489920 4004
rect 489972 3992 489978 4004
rect 491110 3992 491116 4004
rect 489972 3964 491116 3992
rect 489972 3952 489978 3964
rect 491110 3952 491116 3964
rect 491168 3952 491174 4004
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 46716 3896 113174 3924
rect 46716 3884 46722 3896
rect 31294 3816 31300 3868
rect 31352 3856 31358 3868
rect 39298 3856 39304 3868
rect 31352 3828 39304 3856
rect 31352 3816 31358 3828
rect 39298 3816 39304 3828
rect 39356 3816 39362 3868
rect 43070 3816 43076 3868
rect 43128 3856 43134 3868
rect 111978 3856 111984 3868
rect 43128 3828 111984 3856
rect 43128 3816 43134 3828
rect 111978 3816 111984 3828
rect 112036 3816 112042 3868
rect 23014 3748 23020 3800
rect 23072 3788 23078 3800
rect 35158 3788 35164 3800
rect 23072 3760 35164 3788
rect 23072 3748 23078 3760
rect 35158 3748 35164 3760
rect 35216 3748 35222 3800
rect 39574 3748 39580 3800
rect 39632 3788 39638 3800
rect 111886 3788 111892 3800
rect 39632 3760 111892 3788
rect 39632 3748 39638 3760
rect 111886 3748 111892 3760
rect 111944 3748 111950 3800
rect 16853 3723 16911 3729
rect 16853 3689 16865 3723
rect 16899 3720 16911 3723
rect 25498 3720 25504 3732
rect 16899 3692 25504 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 25498 3680 25504 3692
rect 25556 3680 25562 3732
rect 38378 3680 38384 3732
rect 38436 3720 38442 3732
rect 43438 3720 43444 3732
rect 38436 3692 43444 3720
rect 38436 3680 38442 3692
rect 43438 3680 43444 3692
rect 43496 3680 43502 3732
rect 43533 3723 43591 3729
rect 43533 3689 43545 3723
rect 43579 3720 43591 3723
rect 110598 3720 110604 3732
rect 43579 3692 110604 3720
rect 43579 3689 43591 3692
rect 43533 3683 43591 3689
rect 110598 3680 110604 3692
rect 110656 3680 110662 3732
rect 15930 3612 15936 3664
rect 15988 3652 15994 3664
rect 21358 3652 21364 3664
rect 15988 3624 21364 3652
rect 15988 3612 15994 3624
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 32306 3652 32312 3664
rect 26206 3624 32312 3652
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 11698 3584 11704 3596
rect 6512 3556 11704 3584
rect 6512 3544 6518 3556
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 16853 3587 16911 3593
rect 16853 3584 16865 3587
rect 13596 3556 16865 3584
rect 13596 3544 13602 3556
rect 16853 3553 16865 3556
rect 16899 3553 16911 3587
rect 22738 3584 22744 3596
rect 16853 3547 16911 3553
rect 16960 3556 22744 3584
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 15838 3516 15844 3528
rect 10008 3488 15844 3516
rect 10008 3476 10014 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 16960 3516 16988 3556
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 16546 3488 16988 3516
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 7558 3448 7564 3460
rect 1728 3420 7564 3448
rect 1728 3408 1734 3420
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 8754 3408 8760 3460
rect 8812 3448 8818 3460
rect 16546 3448 16574 3488
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 26206 3516 26234 3624
rect 32306 3612 32312 3624
rect 32364 3612 32370 3664
rect 32398 3612 32404 3664
rect 32456 3652 32462 3664
rect 110506 3652 110512 3664
rect 32456 3624 110512 3652
rect 32456 3612 32462 3624
rect 110506 3612 110512 3624
rect 110564 3612 110570 3664
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 109126 3584 109132 3596
rect 28960 3556 109132 3584
rect 28960 3544 28966 3556
rect 109126 3544 109132 3556
rect 109184 3544 109190 3596
rect 18288 3488 26234 3516
rect 18288 3476 18294 3488
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
<<<<<<< HEAD
rect 103793 3519 103851 3525
rect 103793 3516 103805 3519
rect 34532 3488 103805 3516
=======
rect 106829 3519 106887 3525
rect 106829 3516 106841 3519
rect 34532 3488 106841 3516
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 8812 3420 16574 3448
rect 8812 3408 8818 3420
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 34532 3448 34560 3488
<<<<<<< HEAD
rect 103793 3485 103805 3488
rect 103839 3485 103851 3519
rect 105633 3519 105691 3525
rect 105633 3516 105645 3519
rect 103793 3479 103851 3485
rect 103900 3488 105645 3516
rect 103900 3448 103928 3488
rect 105633 3485 105645 3488
rect 105679 3485 105691 3519
rect 105633 3479 105691 3485
=======
rect 106829 3485 106841 3488
rect 106875 3485 106887 3519
rect 106829 3479 106887 3485
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
<<<<<<< HEAD
=======
rect 107657 3519 107715 3525
rect 107657 3485 107669 3519
rect 107703 3516 107715 3519
rect 109218 3516 109224 3528
rect 107703 3488 109224 3516
rect 107703 3485 107715 3488
rect 107657 3479 107715 3485
rect 109218 3476 109224 3488
rect 109276 3476 109282 3528
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111702 3516 111708 3528
rect 110564 3488 111708 3516
rect 110564 3476 110570 3488
rect 111702 3476 111708 3488
rect 111760 3476 111766 3528
rect 113146 3516 113174 3896
rect 140590 3884 140596 3936
rect 140648 3924 140654 3936
rect 157794 3924 157800 3936
rect 140648 3896 157800 3924
rect 140648 3884 140654 3896
rect 157794 3884 157800 3896
rect 157852 3884 157858 3936
rect 158898 3884 158904 3936
rect 158956 3924 158962 3936
rect 177298 3924 177304 3936
rect 158956 3896 177304 3924
rect 158956 3884 158962 3896
rect 177298 3884 177304 3896
rect 177356 3884 177362 3936
rect 192018 3884 192024 3936
rect 192076 3924 192082 3936
rect 206370 3924 206376 3936
rect 192076 3896 206376 3924
rect 192076 3884 192082 3896
rect 206370 3884 206376 3896
rect 206428 3884 206434 3936
rect 209774 3884 209780 3936
rect 209832 3924 209838 3936
rect 209832 3896 224540 3924
rect 209832 3884 209838 3896
rect 131758 3816 131764 3868
rect 131816 3856 131822 3868
rect 162118 3856 162124 3868
rect 131816 3828 162124 3856
rect 131816 3816 131822 3828
rect 162118 3816 162124 3828
rect 162176 3816 162182 3868
rect 170766 3816 170772 3868
rect 170824 3856 170830 3868
rect 178678 3856 178684 3868
rect 170824 3828 178684 3856
rect 170824 3816 170830 3828
rect 178678 3816 178684 3828
rect 178736 3816 178742 3868
rect 184934 3816 184940 3868
rect 184992 3856 184998 3868
rect 196618 3856 196624 3868
rect 184992 3828 196624 3856
rect 184992 3816 184998 3828
rect 196618 3816 196624 3828
rect 196676 3816 196682 3868
rect 206186 3816 206192 3868
rect 206244 3856 206250 3868
rect 224402 3856 224408 3868
rect 206244 3828 224408 3856
rect 206244 3816 206250 3828
rect 224402 3816 224408 3828
rect 224460 3816 224466 3868
rect 224512 3856 224540 3896
rect 227530 3884 227536 3936
rect 227588 3924 227594 3936
rect 231210 3924 231216 3936
rect 227588 3896 231216 3924
rect 227588 3884 227594 3896
rect 231210 3884 231216 3896
rect 231268 3884 231274 3936
rect 255866 3884 255872 3936
rect 255924 3924 255930 3936
rect 336826 3924 336832 3936
rect 255924 3896 336832 3924
rect 255924 3884 255930 3896
rect 336826 3884 336832 3896
rect 336884 3884 336890 3936
<<<<<<< HEAD
=======
rect 352006 3924 352012 3936
rect 345676 3896 352012 3924
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 228450 3856 228456 3868
rect 224512 3828 228456 3856
rect 228450 3816 228456 3828
rect 228508 3816 228514 3868
rect 252370 3816 252376 3868
rect 252428 3856 252434 3868
rect 336734 3856 336740 3868
rect 252428 3828 336740 3856
rect 252428 3816 252434 3828
rect 336734 3816 336740 3828
rect 336792 3816 336798 3868
rect 337289 3859 337347 3865
rect 337289 3825 337301 3859
rect 337335 3856 337347 3859
<<<<<<< HEAD
rect 341150 3856 341156 3868
rect 337335 3828 341156 3856
rect 337335 3825 337347 3828
rect 337289 3819 337347 3825
rect 341150 3816 341156 3828
rect 341208 3816 341214 3868
=======
rect 340966 3856 340972 3868
rect 337335 3828 340972 3856
rect 337335 3825 337347 3828
rect 337289 3819 337347 3825
rect 340966 3816 340972 3828
rect 341024 3816 341030 3868
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 135254 3748 135260 3800
rect 135312 3788 135318 3800
rect 173250 3788 173256 3800
rect 135312 3760 173256 3788
rect 135312 3748 135318 3760
rect 173250 3748 173256 3760
rect 173308 3748 173314 3800
rect 177942 3748 177948 3800
rect 178000 3788 178006 3800
rect 195330 3788 195336 3800
rect 178000 3760 195336 3788
rect 178000 3748 178006 3760
rect 195330 3748 195336 3760
rect 195388 3748 195394 3800
rect 199102 3748 199108 3800
rect 199160 3788 199166 3800
rect 209038 3788 209044 3800
rect 199160 3760 209044 3788
rect 199160 3748 199166 3760
rect 209038 3748 209044 3760
rect 209096 3748 209102 3800
rect 213362 3748 213368 3800
rect 213420 3788 213426 3800
rect 232590 3788 232596 3800
rect 213420 3760 232596 3788
rect 213420 3748 213426 3760
rect 232590 3748 232596 3760
rect 232648 3748 232654 3800
rect 238110 3748 238116 3800
rect 238168 3788 238174 3800
rect 242250 3788 242256 3800
rect 238168 3760 242256 3788
rect 238168 3748 238174 3760
rect 242250 3748 242256 3760
rect 242308 3748 242314 3800
rect 248782 3748 248788 3800
rect 248840 3788 248846 3800
rect 335446 3788 335452 3800
rect 248840 3760 335452 3788
rect 248840 3748 248846 3760
rect 335446 3748 335452 3760
rect 335504 3748 335510 3800
<<<<<<< HEAD
rect 340966 3748 340972 3800
rect 341024 3788 341030 3800
rect 342070 3788 342076 3800
rect 341024 3760 342076 3788
rect 341024 3748 341030 3760
rect 342070 3748 342076 3760
rect 342128 3748 342134 3800
=======
rect 337105 3791 337163 3797
rect 337105 3757 337117 3791
rect 337151 3788 337163 3791
rect 343726 3788 343732 3800
rect 337151 3760 343732 3788
rect 337151 3757 337163 3760
rect 337105 3751 337163 3757
rect 343726 3748 343732 3760
rect 343784 3748 343790 3800
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 142062 3680 142068 3732
rect 142120 3720 142126 3732
rect 160005 3723 160063 3729
rect 160005 3720 160017 3723
rect 142120 3692 160017 3720
rect 142120 3680 142126 3692
rect 160005 3689 160017 3692
rect 160051 3689 160063 3723
rect 160005 3683 160063 3689
rect 160094 3680 160100 3732
rect 160152 3720 160158 3732
<<<<<<< HEAD
rect 316037 3723 316095 3729
rect 316037 3720 316049 3723
rect 160152 3692 316049 3720
rect 160152 3680 160158 3692
rect 316037 3689 316049 3692
rect 316083 3689 316095 3723
rect 316037 3683 316095 3689
rect 316126 3680 316132 3732
rect 316184 3720 316190 3732
rect 316402 3720 316408 3732
rect 316184 3692 316408 3720
rect 316184 3680 316190 3692
rect 316402 3680 316408 3692
rect 316460 3680 316466 3732
rect 333882 3680 333888 3732
rect 333940 3720 333946 3732
rect 345676 3720 345704 3964
rect 352006 3952 352012 3964
rect 352064 3952 352070 4004
rect 361482 3952 361488 4004
rect 361540 3992 361546 4004
rect 376478 3992 376484 4004
rect 361540 3964 376484 3992
rect 361540 3952 361546 3964
rect 376478 3952 376484 3964
rect 376536 3952 376542 4004
rect 382182 3952 382188 4004
rect 382240 3992 382246 4004
rect 479334 3992 479340 4004
rect 382240 3964 479340 3992
rect 382240 3952 382246 3964
rect 479334 3952 479340 3964
rect 479392 3952 479398 4004
rect 349430 3924 349436 3936
rect 349391 3896 349436 3924
rect 349430 3884 349436 3896
rect 349488 3884 349494 3936
=======
rect 318886 3720 318892 3732
rect 160152 3692 318892 3720
rect 160152 3680 160158 3692
rect 318886 3680 318892 3692
rect 318944 3680 318950 3732
rect 333882 3680 333888 3732
rect 333940 3720 333946 3732
rect 345676 3720 345704 3896
rect 352006 3884 352012 3896
rect 352064 3884 352070 3936
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 360838 3884 360844 3936
rect 360896 3924 360902 3936
rect 364610 3924 364616 3936
rect 360896 3896 364616 3924
rect 360896 3884 360902 3896
rect 364610 3884 364616 3896
rect 364668 3884 364674 3936
rect 397362 3884 397368 3936
rect 397420 3924 397426 3936
rect 400309 3927 400367 3933
rect 400309 3924 400321 3927
rect 397420 3896 400321 3924
rect 397420 3884 397426 3896
rect 400309 3893 400321 3896
rect 400355 3893 400367 3927
rect 400309 3887 400367 3893
rect 400401 3927 400459 3933
rect 400401 3893 400413 3927
rect 400447 3924 400459 3927
rect 550266 3924 550272 3936
rect 400447 3896 550272 3924
rect 400447 3893 400459 3896
rect 400401 3887 400459 3893
rect 550266 3884 550272 3896
rect 550324 3884 550330 3936
rect 362862 3816 362868 3868
rect 362920 3856 362926 3868
rect 379974 3856 379980 3868
rect 362920 3828 379980 3856
rect 362920 3816 362926 3828
rect 379974 3816 379980 3828
rect 380032 3816 380038 3868
rect 397270 3816 397276 3868
rect 397328 3856 397334 3868
rect 553762 3856 553768 3868
rect 397328 3828 553768 3856
rect 397328 3816 397334 3828
rect 553762 3816 553768 3828
rect 553820 3816 553826 3868
rect 351914 3788 351920 3800
rect 333940 3692 345704 3720
rect 345768 3760 351920 3788
rect 333940 3680 333946 3692
<<<<<<< HEAD
rect 139210 3612 139216 3664
rect 139268 3652 139274 3664
rect 139268 3624 140176 3652
rect 139268 3612 139274 3624
rect 137830 3544 137836 3596
rect 137888 3584 137894 3596
rect 140038 3584 140044 3596
rect 137888 3556 140044 3584
rect 137888 3544 137894 3556
rect 140038 3544 140044 3556
rect 140096 3544 140102 3596
rect 140148 3584 140176 3624
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 140682 3612 140688 3664
rect 140740 3652 140746 3664
rect 154206 3652 154212 3664
rect 140740 3624 154212 3652
rect 140740 3612 140746 3624
rect 154206 3612 154212 3624
rect 154264 3612 154270 3664
rect 156598 3612 156604 3664
rect 156656 3652 156662 3664
rect 311345 3655 311403 3661
rect 156656 3624 311296 3652
rect 156656 3612 156662 3624
<<<<<<< HEAD
rect 150618 3584 150624 3596
rect 140148 3556 150624 3584
=======
rect 139210 3544 139216 3596
rect 139268 3584 139274 3596
rect 150618 3584 150624 3596
rect 139268 3556 150624 3584
rect 139268 3544 139274 3556
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 150618 3544 150624 3556
rect 150676 3544 150682 3596
rect 153010 3544 153016 3596
rect 153068 3584 153074 3596
rect 311161 3587 311219 3593
rect 311161 3584 311173 3587
rect 153068 3556 311173 3584
rect 153068 3544 153074 3556
rect 311161 3553 311173 3556
rect 311207 3553 311219 3587
rect 311268 3584 311296 3624
rect 311345 3621 311357 3655
rect 311391 3652 311403 3655
rect 317506 3652 317512 3664
rect 311391 3624 317512 3652
rect 311391 3621 311403 3624
rect 311345 3615 311403 3621
rect 317506 3612 317512 3624
rect 317564 3612 317570 3664
rect 319714 3612 319720 3664
rect 319772 3652 319778 3664
rect 319772 3624 325694 3652
rect 319772 3612 319778 3624
rect 312541 3587 312599 3593
rect 312541 3584 312553 3587
rect 311268 3556 312553 3584
rect 311161 3547 311219 3553
rect 312541 3553 312553 3556
rect 312587 3553 312599 3587
rect 312541 3547 312599 3553
rect 312630 3544 312636 3596
rect 312688 3584 312694 3596
rect 313182 3584 313188 3596
rect 312688 3556 313188 3584
rect 312688 3544 312694 3556
rect 313182 3544 313188 3556
rect 313240 3544 313246 3596
rect 313277 3587 313335 3593
rect 313277 3553 313289 3587
rect 313323 3584 313335 3587
rect 316129 3587 316187 3593
rect 316129 3584 316141 3587
rect 313323 3556 316141 3584
rect 313323 3553 313335 3556
rect 313277 3547 313335 3553
rect 316129 3553 316141 3556
rect 316175 3553 316187 3587
rect 316129 3547 316187 3553
rect 316218 3544 316224 3596
rect 316276 3584 316282 3596
<<<<<<< HEAD
rect 316276 3556 324452 3584
=======
rect 316276 3556 317736 3584
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 316276 3544 316282 3556
rect 113266 3516 113272 3528
rect 113146 3488 113272 3516
rect 113266 3476 113272 3488
rect 113324 3476 113330 3528
<<<<<<< HEAD
rect 113821 3519 113879 3525
rect 113821 3485 113833 3519
rect 113867 3516 113879 3519
rect 118970 3516 118976 3528
rect 113867 3488 118976 3516
rect 113867 3485 113879 3488
rect 113821 3479 113879 3485
rect 118970 3476 118976 3488
rect 119028 3476 119034 3528
=======
rect 114002 3476 114008 3528
rect 114060 3516 114066 3528
rect 114462 3516 114468 3528
rect 114060 3488 114468 3516
rect 114060 3476 114066 3488
rect 114462 3476 114468 3488
rect 114520 3476 114526 3528
rect 116397 3519 116455 3525
rect 116397 3485 116409 3519
rect 116443 3516 116455 3519
rect 121638 3516 121644 3528
rect 116443 3488 121644 3516
rect 116443 3485 116455 3488
rect 116397 3479 116455 3485
rect 121638 3476 121644 3488
rect 121696 3476 121702 3528
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 126882 3516 126888 3528
rect 125928 3488 126888 3516
rect 125928 3476 125934 3488
rect 126882 3476 126888 3488
rect 126940 3476 126946 3528
<<<<<<< HEAD
=======
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 129550 3516 129556 3528
rect 127032 3488 129556 3516
rect 127032 3476 127038 3488
rect 129550 3476 129556 3488
rect 129608 3476 129614 3528
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 130562 3476 130568 3528
rect 130620 3516 130626 3528
rect 131022 3516 131028 3528
rect 130620 3488 131028 3516
rect 130620 3476 130626 3488
rect 131022 3476 131028 3488
rect 131080 3476 131086 3528
rect 132954 3476 132960 3528
rect 133012 3516 133018 3528
rect 133782 3516 133788 3528
rect 133012 3488 133788 3516
rect 133012 3476 133018 3488
rect 133782 3476 133788 3488
rect 133840 3476 133846 3528
<<<<<<< HEAD
rect 134518 3516 134524 3528
rect 133892 3488 134524 3516
rect 24268 3420 34560 3448
rect 35866 3420 103928 3448
rect 103977 3451 104035 3457
rect 24268 3408 24274 3420
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 35866 3380 35894 3420
rect 103977 3417 103989 3451
rect 104023 3448 104035 3451
rect 114554 3448 114560 3460
rect 104023 3420 114560 3448
rect 104023 3417 104035 3420
rect 103977 3411 104035 3417
rect 114554 3408 114560 3420
rect 114612 3408 114618 3460
rect 116397 3451 116455 3457
rect 116397 3417 116409 3451
rect 116443 3448 116455 3451
rect 121638 3448 121644 3460
rect 116443 3420 121644 3448
rect 116443 3417 116455 3420
rect 116397 3411 116455 3417
rect 121638 3408 121644 3420
rect 121696 3408 121702 3460
rect 128170 3408 128176 3460
rect 128228 3448 128234 3460
rect 133892 3448 133920 3488
rect 134518 3476 134524 3488
rect 134576 3476 134582 3528
rect 139302 3476 139308 3528
rect 139360 3516 139366 3528
rect 147122 3516 147128 3528
rect 139360 3488 147128 3516
rect 139360 3476 139366 3488
rect 147122 3476 147128 3488
rect 147180 3476 147186 3528
=======
rect 141234 3476 141240 3528
rect 141292 3516 141298 3528
rect 141970 3516 141976 3528
rect 141292 3488 141976 3516
rect 141292 3476 141298 3488
rect 141970 3476 141976 3488
rect 142028 3476 142034 3528
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148962 3516 148968 3528
rect 148376 3488 148968 3516
rect 148376 3476 148382 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 149514 3476 149520 3528
rect 149572 3516 149578 3528
<<<<<<< HEAD
rect 316313 3519 316371 3525
rect 149572 3488 316172 3516
rect 149572 3476 149578 3488
rect 316144 3460 316172 3488
rect 316313 3485 316325 3519
rect 316359 3516 316371 3519
rect 317598 3516 317604 3528
rect 316359 3488 317604 3516
rect 316359 3485 316371 3488
rect 316313 3479 316371 3485
rect 317598 3476 317604 3488
rect 317656 3476 317662 3528
rect 128228 3420 133920 3448
rect 128228 3408 128234 3420
rect 134150 3408 134156 3460
rect 134208 3448 134214 3460
rect 135162 3448 135168 3460
rect 134208 3420 135168 3448
rect 134208 3408 134214 3420
rect 135162 3408 135168 3420
rect 135220 3408 135226 3460
=======
rect 316402 3516 316408 3528
rect 149572 3488 316408 3516
rect 149572 3476 149578 3488
rect 316402 3476 316408 3488
rect 316460 3476 316466 3528
rect 107838 3448 107844 3460
rect 24268 3420 34560 3448
rect 35866 3420 107844 3448
rect 24268 3408 24274 3420
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 35866 3380 35894 3420
rect 107838 3408 107844 3420
rect 107896 3408 107902 3460
rect 108301 3451 108359 3457
rect 108301 3417 108313 3451
rect 108347 3448 108359 3451
rect 114554 3448 114560 3460
rect 108347 3420 114560 3448
rect 108347 3417 108359 3420
rect 108301 3411 108359 3417
rect 114554 3408 114560 3420
rect 114612 3408 114618 3460
rect 116581 3451 116639 3457
rect 116581 3417 116593 3451
rect 116627 3448 116639 3451
rect 121546 3448 121552 3460
rect 116627 3420 121552 3448
rect 116627 3417 116639 3420
rect 116581 3411 116639 3417
rect 121546 3408 121552 3420
rect 121604 3408 121610 3460
rect 128170 3408 128176 3460
rect 128228 3448 128234 3460
rect 134518 3448 134524 3460
rect 128228 3420 134524 3448
rect 128228 3408 128234 3420
rect 134518 3408 134524 3420
rect 134576 3408 134582 3460
rect 139302 3408 139308 3460
rect 139360 3448 139366 3460
rect 139360 3420 142154 3448
rect 139360 3408 139366 3420
rect 19484 3352 35894 3380
rect 19484 3340 19490 3352
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 50154 3340 50160 3392
rect 50212 3380 50218 3392
rect 50982 3380 50988 3392
rect 50212 3352 50988 3380
rect 50212 3340 50218 3352
rect 50982 3340 50988 3352
rect 51040 3340 51046 3392
rect 67910 3340 67916 3392
rect 67968 3380 67974 3392
rect 117406 3380 117412 3392
rect 67968 3352 117412 3380
rect 67968 3340 67974 3352
rect 117406 3340 117412 3352
rect 117464 3340 117470 3392
rect 137830 3340 137836 3392
rect 137888 3380 137894 3392
rect 140038 3380 140044 3392
rect 137888 3352 140044 3380
rect 137888 3340 137894 3352
rect 140038 3340 140044 3352
rect 140096 3340 140102 3392
rect 142126 3380 142154 3420
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 145926 3408 145932 3460
rect 145984 3448 145990 3460
rect 316034 3448 316040 3460
rect 145984 3420 316040 3448
rect 145984 3408 145990 3420
rect 316034 3408 316040 3420
rect 316092 3408 316098 3460
<<<<<<< HEAD
rect 316126 3408 316132 3460
rect 316184 3408 316190 3460
rect 316221 3451 316279 3457
rect 316221 3417 316233 3451
rect 316267 3448 316279 3451
rect 318886 3448 318892 3460
rect 316267 3420 318892 3448
rect 316267 3417 316279 3420
rect 316221 3411 316279 3417
rect 318886 3408 318892 3420
rect 318944 3408 318950 3460
rect 323302 3408 323308 3460
rect 323360 3448 323366 3460
rect 324222 3448 324228 3460
rect 323360 3420 324228 3448
rect 323360 3408 323366 3420
rect 324222 3408 324228 3420
rect 324280 3408 324286 3460
rect 324424 3448 324452 3556
=======
rect 316129 3451 316187 3457
rect 316129 3417 316141 3451
rect 316175 3448 316187 3451
rect 317598 3448 317604 3460
rect 316175 3420 317604 3448
rect 316175 3417 316187 3420
rect 316129 3411 316187 3417
rect 317598 3408 317604 3420
rect 317656 3408 317662 3460
rect 317708 3448 317736 3556
rect 323302 3476 323308 3528
rect 323360 3516 323366 3528
rect 324222 3516 324228 3528
rect 323360 3488 324228 3516
rect 323360 3476 323366 3488
rect 324222 3476 324228 3488
rect 324280 3476 324286 3528
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 325666 3516 325694 3624
rect 330386 3612 330392 3664
rect 330444 3652 330450 3664
rect 345768 3652 345796 3760
rect 351914 3748 351920 3760
rect 351972 3748 351978 3800
rect 362770 3748 362776 3800
rect 362828 3788 362834 3800
rect 383562 3788 383568 3800
rect 362828 3760 383568 3788
rect 362828 3748 362834 3760
rect 383562 3748 383568 3760
rect 383620 3748 383626 3800
rect 395982 3748 395988 3800
rect 396040 3788 396046 3800
rect 399849 3791 399907 3797
rect 399849 3788 399861 3791
rect 396040 3760 399861 3788
rect 396040 3748 396046 3760
rect 399849 3757 399861 3760
rect 399895 3757 399907 3791
rect 399849 3751 399907 3757
rect 399938 3748 399944 3800
rect 399996 3788 400002 3800
rect 400217 3791 400275 3797
rect 400217 3788 400229 3791
rect 399996 3760 400229 3788
rect 399996 3748 400002 3760
rect 400217 3757 400229 3760
rect 400263 3757 400275 3791
rect 400217 3751 400275 3757
rect 400309 3791 400367 3797
rect 400309 3757 400321 3791
rect 400355 3788 400367 3791
rect 557350 3788 557356 3800
rect 400355 3760 557356 3788
rect 400355 3757 400367 3760
rect 400309 3751 400367 3757
rect 557350 3748 557356 3760
rect 557408 3748 557414 3800
rect 364242 3680 364248 3732
rect 364300 3720 364306 3732
rect 387150 3720 387156 3732
rect 364300 3692 387156 3720
rect 364300 3680 364306 3692
rect 387150 3680 387156 3692
rect 387208 3680 387214 3732
rect 398742 3680 398748 3732
rect 398800 3720 398806 3732
rect 560846 3720 560852 3732
rect 398800 3692 560852 3720
rect 398800 3680 398806 3692
rect 560846 3680 560852 3692
rect 560904 3680 560910 3732
rect 350718 3652 350724 3664
rect 330444 3624 345796 3652
rect 345860 3624 350724 3652
rect 330444 3612 330450 3624
rect 326798 3544 326804 3596
rect 326856 3584 326862 3596
rect 345860 3584 345888 3624
rect 350718 3612 350724 3624
rect 350776 3612 350782 3664
rect 353938 3612 353944 3664
rect 353996 3652 354002 3664
rect 357526 3652 357532 3664
rect 353996 3624 357532 3652
rect 353996 3612 354002 3624
rect 357526 3612 357532 3624
rect 357584 3612 357590 3664
rect 360010 3612 360016 3664
rect 360068 3652 360074 3664
rect 360068 3624 362448 3652
rect 360068 3612 360074 3624
rect 326856 3556 345888 3584
rect 326856 3544 326862 3556
rect 348050 3544 348056 3596
rect 348108 3584 348114 3596
rect 354766 3584 354772 3596
rect 348108 3556 354772 3584
rect 348108 3544 348114 3556
rect 354766 3544 354772 3556
rect 354824 3544 354830 3596
rect 358630 3544 358636 3596
rect 358688 3584 358694 3596
rect 362310 3584 362316 3596
rect 358688 3556 362316 3584
rect 358688 3544 358694 3556
rect 362310 3544 362316 3556
rect 362368 3544 362374 3596
rect 362420 3584 362448 3624
rect 364150 3612 364156 3664
rect 364208 3652 364214 3664
rect 390646 3652 390652 3664
rect 364208 3624 390652 3652
rect 364208 3612 364214 3624
rect 390646 3612 390652 3624
rect 390704 3612 390710 3664
rect 398650 3612 398656 3664
rect 398708 3652 398714 3664
rect 564434 3652 564440 3664
rect 398708 3624 564440 3652
rect 398708 3612 398714 3624
rect 564434 3612 564440 3624
rect 564492 3612 564498 3664
rect 369394 3584 369400 3596
rect 362420 3556 369400 3584
rect 369394 3544 369400 3556
rect 369452 3544 369458 3596
rect 394234 3584 394240 3596
rect 369504 3556 394240 3584
rect 349154 3516 349160 3528
rect 325666 3488 349160 3516
rect 349154 3476 349160 3488
rect 349212 3476 349218 3528
rect 355226 3476 355232 3528
rect 355284 3516 355290 3528
rect 356238 3516 356244 3528
rect 355284 3488 356244 3516
rect 355284 3476 355290 3488
rect 356238 3476 356244 3488
rect 356296 3476 356302 3528
rect 357434 3476 357440 3528
rect 357492 3516 357498 3528
rect 358722 3516 358728 3528
rect 357492 3488 358728 3516
rect 357492 3476 357498 3488
rect 358722 3476 358728 3488
rect 358780 3476 358786 3528
rect 365622 3476 365628 3528
rect 365680 3516 365686 3528
rect 369504 3516 369532 3556
rect 394234 3544 394240 3556
rect 394292 3544 394298 3596
rect 400030 3544 400036 3596
rect 400088 3584 400094 3596
rect 568022 3584 568028 3596
rect 400088 3556 568028 3584
rect 400088 3544 400094 3556
rect 568022 3544 568028 3556
rect 568080 3544 568086 3596
rect 397730 3516 397736 3528
rect 365680 3488 369532 3516
rect 369596 3488 397736 3516
rect 365680 3476 365686 3488
<<<<<<< HEAD
rect 349433 3451 349491 3457
rect 349433 3448 349445 3451
rect 324424 3420 349445 3448
rect 349433 3417 349445 3420
rect 349479 3417 349491 3451
rect 349433 3411 349491 3417
=======
rect 349430 3448 349436 3460
rect 317708 3420 349436 3448
rect 349430 3408 349436 3420
rect 349488 3408 349494 3460
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 354122 3408 354128 3460
rect 354180 3448 354186 3460
rect 361114 3448 361120 3460
rect 354180 3420 361120 3448
rect 354180 3408 354186 3420
rect 361114 3408 361120 3420
rect 361172 3408 361178 3460
rect 365530 3408 365536 3460
rect 365588 3448 365594 3460
rect 369596 3448 369624 3488
rect 397730 3476 397736 3488
rect 397788 3476 397794 3528
rect 398834 3476 398840 3528
rect 398892 3516 398898 3528
rect 400122 3516 400128 3528
rect 398892 3488 400128 3516
rect 398892 3476 398898 3488
rect 400122 3476 400128 3488
rect 400180 3476 400186 3528
rect 400217 3519 400275 3525
rect 400217 3485 400229 3519
rect 400263 3516 400275 3519
rect 571518 3516 571524 3528
rect 400263 3488 571524 3516
rect 400263 3485 400275 3488
rect 400217 3479 400275 3485
rect 571518 3476 571524 3488
rect 571576 3476 571582 3528
rect 401318 3448 401324 3460
rect 365588 3420 369624 3448
rect 373966 3420 401324 3448
rect 365588 3408 365594 3420
<<<<<<< HEAD
rect 19484 3352 35894 3380
rect 19484 3340 19490 3352
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 50154 3340 50160 3392
rect 50212 3380 50218 3392
rect 50982 3380 50988 3392
rect 50212 3352 50988 3380
rect 50212 3340 50218 3352
rect 50982 3340 50988 3352
rect 51040 3340 51046 3392
rect 72602 3340 72608 3392
rect 72660 3380 72666 3392
rect 73062 3380 73068 3392
rect 72660 3352 73068 3380
rect 72660 3340 72666 3352
rect 73062 3340 73068 3352
rect 73120 3340 73126 3392
rect 117406 3380 117412 3392
rect 73264 3352 117412 3380
rect 35986 3272 35992 3324
rect 36044 3312 36050 3324
rect 43533 3315 43591 3321
rect 43533 3312 43545 3315
rect 36044 3284 43545 3312
rect 36044 3272 36050 3284
rect 43533 3281 43545 3284
rect 43579 3281 43591 3315
rect 43533 3275 43591 3281
rect 67910 3204 67916 3256
rect 67968 3244 67974 3256
rect 73264 3244 73292 3352
rect 117406 3340 117412 3352
rect 117464 3340 117470 3392
=======
rect 147122 3380 147128 3392
rect 142126 3352 147128 3380
rect 147122 3340 147128 3352
rect 147180 3340 147186 3392
rect 155402 3340 155408 3392
rect 155460 3380 155466 3392
rect 155862 3380 155868 3392
rect 155460 3352 155868 3380
rect 155460 3340 155466 3352
rect 155862 3340 155868 3352
rect 155920 3340 155926 3392
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 160005 3383 160063 3389
rect 160005 3349 160017 3383
rect 160051 3380 160063 3383
rect 161290 3380 161296 3392
rect 160051 3352 161296 3380
rect 160051 3349 160063 3352
rect 160005 3343 160063 3349
rect 161290 3340 161296 3352
rect 161348 3340 161354 3392
rect 163682 3340 163688 3392
rect 163740 3380 163746 3392
rect 164142 3380 164148 3392
rect 163740 3352 164148 3380
rect 163740 3340 163746 3352
rect 164142 3340 164148 3352
rect 164200 3340 164206 3392
rect 173158 3340 173164 3392
rect 173216 3380 173222 3392
rect 173618 3380 173624 3392
rect 173216 3352 173624 3380
rect 173216 3340 173222 3352
rect 173618 3340 173624 3352
rect 173676 3340 173682 3392
rect 174262 3340 174268 3392
rect 174320 3380 174326 3392
rect 175090 3380 175096 3392
rect 174320 3352 175096 3380
rect 174320 3340 174326 3352
rect 175090 3340 175096 3352
rect 175148 3340 175154 3392
rect 176654 3340 176660 3392
rect 176712 3380 176718 3392
rect 177850 3380 177856 3392
rect 176712 3352 177856 3380
rect 176712 3340 176718 3352
rect 177850 3340 177856 3352
rect 177908 3340 177914 3392
rect 181438 3340 181444 3392
rect 181496 3380 181502 3392
rect 181898 3380 181904 3392
rect 181496 3352 181904 3380
rect 181496 3340 181502 3352
rect 181898 3340 181904 3352
rect 181956 3340 181962 3392
<<<<<<< HEAD
=======
rect 190822 3340 190828 3392
rect 190880 3380 190886 3392
rect 191558 3380 191564 3392
rect 190880 3352 191564 3380
rect 190880 3340 190886 3352
rect 191558 3340 191564 3352
rect 191616 3340 191622 3392
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 197906 3340 197912 3392
rect 197964 3380 197970 3392
rect 198550 3380 198556 3392
rect 197964 3352 198556 3380
rect 197964 3340 197970 3352
rect 198550 3340 198556 3352
rect 198608 3340 198614 3392
<<<<<<< HEAD
=======
rect 201494 3340 201500 3392
rect 201552 3380 201558 3392
rect 202506 3380 202512 3392
rect 201552 3352 202512 3380
rect 201552 3340 201558 3352
rect 202506 3340 202512 3352
rect 202564 3340 202570 3392
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 208578 3340 208584 3392
rect 208636 3380 208642 3392
rect 209682 3380 209688 3392
rect 208636 3352 209688 3380
rect 208636 3340 208642 3352
rect 209682 3340 209688 3352
rect 209740 3340 209746 3392
rect 226334 3340 226340 3392
rect 226392 3380 226398 3392
rect 227622 3380 227628 3392
rect 226392 3352 227628 3380
rect 226392 3340 226398 3352
rect 227622 3340 227628 3352
rect 227680 3340 227686 3392
rect 231026 3340 231032 3392
rect 231084 3380 231090 3392
rect 231762 3380 231768 3392
rect 231084 3352 231768 3380
rect 231084 3340 231090 3352
rect 231762 3340 231768 3352
rect 231820 3340 231826 3392
rect 233418 3340 233424 3392
rect 233476 3380 233482 3392
rect 234522 3380 234528 3392
rect 233476 3352 234528 3380
rect 233476 3340 233482 3352
rect 234522 3340 234528 3352
rect 234580 3340 234586 3392
<<<<<<< HEAD
rect 259454 3340 259460 3392
rect 259512 3380 259518 3392
rect 260650 3380 260656 3392
rect 259512 3352 260656 3380
rect 259512 3340 259518 3352
rect 260650 3340 260656 3352
rect 260708 3340 260714 3392
rect 270034 3340 270040 3392
rect 270092 3380 270098 3392
rect 270092 3352 337424 3380
rect 270092 3340 270098 3352
rect 67968 3216 73292 3244
rect 74506 3284 113956 3312
rect 67968 3204 67974 3216
rect 71498 3136 71504 3188
rect 71556 3176 71562 3188
rect 74506 3176 74534 3284
rect 74994 3204 75000 3256
rect 75052 3244 75058 3256
rect 113821 3247 113879 3253
rect 113821 3244 113833 3247
rect 75052 3216 113833 3244
rect 75052 3204 75058 3216
rect 113821 3213 113833 3216
rect 113867 3213 113879 3247
rect 113928 3244 113956 3284
rect 114002 3272 114008 3324
rect 114060 3312 114066 3324
rect 114462 3312 114468 3324
rect 114060 3284 114468 3312
rect 114060 3272 114066 3284
rect 114462 3272 114468 3284
rect 114520 3272 114526 3324
rect 116581 3315 116639 3321
rect 116581 3281 116593 3315
rect 116627 3312 116639 3315
rect 121546 3312 121552 3324
rect 116627 3284 121552 3312
rect 116627 3281 116639 3284
rect 116581 3275 116639 3281
rect 121546 3272 121552 3284
rect 121604 3272 121610 3324
rect 151814 3272 151820 3324
rect 151872 3312 151878 3324
rect 160738 3312 160744 3324
rect 151872 3284 160744 3312
rect 151872 3272 151878 3284
rect 160738 3272 160744 3284
rect 160796 3272 160802 3324
rect 273622 3272 273628 3324
rect 273680 3312 273686 3324
rect 337289 3315 337347 3321
rect 337289 3312 337301 3315
rect 273680 3284 337301 3312
rect 273680 3272 273686 3284
rect 337289 3281 337301 3284
rect 337335 3281 337347 3315
rect 337396 3312 337424 3352
rect 337470 3340 337476 3392
rect 337528 3380 337534 3392
rect 338022 3380 338028 3392
rect 337528 3352 338028 3380
rect 337528 3340 337534 3352
rect 338022 3340 338028 3352
rect 338080 3340 338086 3392
rect 339678 3312 339684 3324
rect 337396 3284 339684 3312
rect 337289 3275 337347 3281
rect 339678 3272 339684 3284
rect 339736 3272 339742 3324
=======
rect 234614 3340 234620 3392
rect 234672 3380 234678 3392
rect 235902 3380 235908 3392
rect 234672 3352 235908 3380
rect 234672 3340 234678 3352
rect 235902 3340 235908 3352
rect 235960 3340 235966 3392
rect 270034 3340 270040 3392
rect 270092 3380 270098 3392
rect 339678 3380 339684 3392
rect 270092 3352 339684 3380
rect 270092 3340 270098 3352
rect 339678 3340 339684 3352
rect 339736 3340 339742 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 342257 3383 342315 3389
rect 342257 3349 342269 3383
rect 342303 3380 342315 3383
rect 346486 3380 346492 3392
rect 342303 3352 346492 3380
rect 342303 3349 342315 3352
rect 342257 3343 342315 3349
rect 346486 3340 346492 3352
rect 346544 3340 346550 3392
rect 35986 3272 35992 3324
rect 36044 3312 36050 3324
rect 43533 3315 43591 3321
rect 43533 3312 43545 3315
rect 36044 3284 43545 3312
rect 36044 3272 36050 3284
rect 43533 3281 43545 3284
rect 43579 3281 43591 3315
rect 43533 3275 43591 3281
rect 71498 3272 71504 3324
rect 71556 3312 71562 3324
rect 117314 3312 117320 3324
rect 71556 3284 117320 3312
rect 71556 3272 71562 3284
rect 117314 3272 117320 3284
rect 117372 3272 117378 3324
rect 273622 3272 273628 3324
rect 273680 3312 273686 3324
rect 273680 3284 337424 3312
rect 273680 3272 273686 3284
rect 72602 3204 72608 3256
rect 72660 3244 72666 3256
rect 73062 3244 73068 3256
rect 72660 3216 73068 3244
rect 72660 3204 72666 3216
rect 73062 3204 73068 3216
rect 73120 3204 73126 3256
rect 74994 3204 75000 3256
rect 75052 3244 75058 3256
rect 118970 3244 118976 3256
rect 75052 3216 118976 3244
rect 75052 3204 75058 3216
rect 118970 3204 118976 3216
rect 119028 3204 119034 3256
rect 277118 3204 277124 3256
rect 277176 3244 277182 3256
rect 337289 3247 337347 3253
rect 337289 3244 337301 3247
rect 277176 3216 337301 3244
rect 277176 3204 277182 3216
rect 337289 3213 337301 3216
rect 337335 3213 337347 3247
rect 337289 3207 337347 3213
rect 41874 3136 41880 3188
rect 41932 3176 41938 3188
rect 42794 3176 42800 3188
rect 41932 3148 42800 3176
rect 41932 3136 41938 3148
rect 42794 3136 42800 3148
rect 42852 3136 42858 3188
rect 78582 3136 78588 3188
rect 78640 3176 78646 3188
rect 118694 3176 118700 3188
rect 78640 3148 118700 3176
rect 78640 3136 78646 3148
rect 118694 3136 118700 3148
rect 118752 3136 118758 3188
rect 134150 3136 134156 3188
rect 134208 3176 134214 3188
rect 135162 3176 135168 3188
rect 134208 3148 135168 3176
rect 134208 3136 134214 3148
rect 135162 3136 135168 3148
rect 135220 3136 135226 3188
rect 166074 3136 166080 3188
rect 166132 3176 166138 3188
rect 170398 3176 170404 3188
rect 166132 3148 170404 3176
rect 166132 3136 166138 3148
rect 170398 3136 170404 3148
rect 170456 3136 170462 3188
rect 284294 3136 284300 3188
rect 284352 3176 284358 3188
rect 337396 3176 337424 3284
rect 337470 3272 337476 3324
rect 337528 3312 337534 3324
rect 338022 3312 338028 3324
rect 337528 3284 338028 3312
rect 337528 3272 337534 3284
rect 338022 3272 338028 3284
rect 338080 3272 338086 3324
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 366818 3272 366824 3324
rect 366876 3312 366882 3324
rect 373966 3312 373994 3420
rect 401318 3408 401324 3420
rect 401376 3408 401382 3460
rect 401502 3408 401508 3460
rect 401560 3448 401566 3460
rect 575106 3448 575112 3460
rect 401560 3420 575112 3448
rect 401560 3408 401566 3420
rect 575106 3408 575112 3420
rect 575164 3408 575170 3460
rect 378042 3340 378048 3392
rect 378100 3380 378106 3392
rect 458082 3380 458088 3392
rect 378100 3352 458088 3380
rect 378100 3340 378106 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
<<<<<<< HEAD
rect 489914 3340 489920 3392
rect 489972 3380 489978 3392
rect 491110 3380 491116 3392
rect 489972 3352 491116 3380
rect 489972 3340 489978 3352
rect 491110 3340 491116 3352
rect 491168 3340 491174 3392
rect 506474 3340 506480 3392
rect 506532 3380 506538 3392
rect 507670 3380 507676 3392
rect 506532 3352 507676 3380
rect 506532 3340 506538 3352
rect 507670 3340 507676 3352
rect 507728 3340 507734 3392
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 530578 3340 530584 3392
rect 530636 3380 530642 3392
rect 532510 3380 532516 3392
rect 530636 3352 532516 3380
rect 530636 3340 530642 3352
rect 532510 3340 532516 3352
rect 532568 3340 532574 3392
rect 366876 3284 373994 3312
rect 366876 3272 366882 3284
rect 375190 3272 375196 3324
rect 375248 3312 375254 3324
rect 375248 3284 375420 3312
rect 375248 3272 375254 3284
<<<<<<< HEAD
rect 117314 3244 117320 3256
rect 113928 3216 117320 3244
rect 113821 3207 113879 3213
rect 117314 3204 117320 3216
rect 117372 3204 117378 3256
rect 277118 3204 277124 3256
rect 277176 3244 277182 3256
rect 340874 3244 340880 3256
rect 277176 3216 340880 3244
rect 277176 3204 277182 3216
rect 340874 3204 340880 3216
rect 340932 3204 340938 3256
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 373994 3204 374000 3256
rect 374052 3244 374058 3256
rect 375282 3244 375288 3256
rect 374052 3216 375288 3244
rect 374052 3204 374058 3216
rect 375282 3204 375288 3216
rect 375340 3204 375346 3256
rect 375392 3244 375420 3284
rect 376662 3272 376668 3324
rect 376720 3312 376726 3324
rect 450906 3312 450912 3324
rect 376720 3284 450912 3312
rect 376720 3272 376726 3284
rect 450906 3272 450912 3284
rect 450964 3272 450970 3324
rect 443822 3244 443828 3256
rect 375392 3216 443828 3244
rect 443822 3204 443828 3216
rect 443880 3204 443886 3256
<<<<<<< HEAD
rect 71556 3148 74534 3176
rect 71556 3136 71562 3148
rect 78582 3136 78588 3188
rect 78640 3176 78646 3188
rect 118694 3176 118700 3188
rect 78640 3148 118700 3176
rect 78640 3136 78646 3148
rect 118694 3136 118700 3148
rect 118752 3136 118758 3188
rect 155402 3136 155408 3188
rect 155460 3176 155466 3188
rect 155862 3176 155868 3188
rect 155460 3148 155868 3176
rect 155460 3136 155466 3148
rect 155862 3136 155868 3148
rect 155920 3136 155926 3188
rect 166074 3136 166080 3188
rect 166132 3176 166138 3188
rect 170398 3176 170404 3188
rect 166132 3148 170404 3176
rect 166132 3136 166138 3148
rect 170398 3136 170404 3148
rect 170456 3136 170462 3188
rect 234614 3136 234620 3188
rect 234672 3176 234678 3188
rect 235902 3176 235908 3188
rect 234672 3148 235908 3176
rect 234672 3136 234678 3148
rect 235902 3136 235908 3148
rect 235960 3136 235966 3188
rect 284294 3136 284300 3188
rect 284352 3176 284358 3188
rect 342438 3176 342444 3188
rect 284352 3148 342444 3176
rect 284352 3136 284358 3148
rect 342438 3136 342444 3148
rect 342496 3136 342502 3188
rect 360102 3136 360108 3188
rect 360160 3176 360166 3188
rect 365806 3176 365812 3188
rect 360160 3148 365812 3176
rect 360160 3136 360166 3148
rect 365806 3136 365812 3148
rect 365864 3136 365870 3188
rect 373902 3136 373908 3188
rect 373960 3176 373966 3188
rect 436738 3176 436744 3188
rect 373960 3148 436744 3176
rect 373960 3136 373966 3148
rect 436738 3136 436744 3148
rect 436796 3136 436802 3188
=======
rect 341150 3176 341156 3188
rect 284352 3148 337332 3176
rect 337396 3148 341156 3176
rect 284352 3136 284358 3148
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 12342 3068 12348 3120
rect 12400 3108 12406 3120
rect 14458 3108 14464 3120
rect 12400 3080 14464 3108
rect 12400 3068 12406 3080
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 82078 3068 82084 3120
rect 82136 3108 82142 3120
rect 120258 3108 120264 3120
rect 82136 3080 120264 3108
rect 82136 3068 82142 3080
rect 120258 3068 120264 3080
rect 120316 3068 120322 3120
<<<<<<< HEAD
rect 126974 3068 126980 3120
rect 127032 3108 127038 3120
rect 129642 3108 129648 3120
rect 127032 3080 129648 3108
rect 127032 3068 127038 3080
rect 129642 3068 129648 3080
rect 129700 3068 129706 3120
rect 201494 3068 201500 3120
rect 201552 3108 201558 3120
rect 202506 3108 202512 3120
rect 201552 3080 202512 3108
rect 201552 3068 201558 3080
rect 202506 3068 202512 3080
rect 202564 3068 202570 3120
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 280706 3068 280712 3120
rect 280764 3108 280770 3120
rect 281442 3108 281448 3120
rect 280764 3080 281448 3108
rect 280764 3068 280770 3080
rect 281442 3068 281448 3080
rect 281500 3068 281506 3120
rect 287790 3068 287796 3120
rect 287848 3108 287854 3120
<<<<<<< HEAD
rect 343634 3108 343640 3120
rect 287848 3080 343640 3108
rect 287848 3068 287854 3080
rect 343634 3068 343640 3080
rect 343692 3068 343698 3120
rect 371142 3068 371148 3120
rect 371200 3108 371206 3120
rect 426158 3108 426164 3120
rect 371200 3080 426164 3108
rect 371200 3068 371206 3080
rect 426158 3068 426164 3080
rect 426216 3068 426222 3120
rect 431954 3068 431960 3120
rect 432012 3108 432018 3120
rect 433242 3108 433248 3120
rect 432012 3080 433248 3108
rect 432012 3068 432018 3080
rect 433242 3068 433248 3080
rect 433300 3068 433306 3120
=======
rect 337304 3108 337332 3148
rect 341150 3136 341156 3148
rect 341208 3136 341214 3188
rect 360102 3136 360108 3188
rect 360160 3176 360166 3188
rect 365806 3176 365812 3188
rect 360160 3148 365812 3176
rect 360160 3136 360166 3148
rect 365806 3136 365812 3148
rect 365864 3136 365870 3188
rect 373902 3136 373908 3188
rect 373960 3176 373966 3188
rect 436738 3176 436744 3188
rect 373960 3148 436744 3176
rect 373960 3136 373966 3148
rect 436738 3136 436744 3148
rect 436796 3136 436802 3188
rect 342438 3108 342444 3120
rect 287848 3080 337240 3108
rect 337304 3080 342444 3108
rect 287848 3068 287854 3080
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 85666 3000 85672 3052
rect 85724 3040 85730 3052
rect 85724 3012 116716 3040
rect 85724 3000 85730 3012
rect 89162 2932 89168 2984
rect 89220 2972 89226 2984
rect 116581 2975 116639 2981
rect 116581 2972 116593 2975
rect 89220 2944 116593 2972
rect 89220 2932 89226 2944
rect 116581 2941 116593 2944
rect 116627 2941 116639 2975
rect 116688 2972 116716 3012
rect 117590 3000 117596 3052
rect 117648 3040 117654 3052
rect 119338 3040 119344 3052
rect 117648 3012 119344 3040
rect 117648 3000 117654 3012
rect 119338 3000 119344 3012
rect 119396 3000 119402 3052
<<<<<<< HEAD
rect 141234 3000 141240 3052
rect 141292 3040 141298 3052
rect 141970 3040 141976 3052
rect 141292 3012 141976 3040
rect 141292 3000 141298 3012
rect 141970 3000 141976 3012
rect 142028 3000 142034 3052
rect 343726 3040 343732 3052
rect 296686 3012 343732 3040
=======
rect 137738 3000 137744 3052
rect 137796 3040 137802 3052
rect 143534 3040 143540 3052
rect 137796 3012 143540 3040
rect 137796 3000 137802 3012
rect 143534 3000 143540 3012
rect 143592 3000 143598 3052
rect 337105 3043 337163 3049
rect 337105 3040 337117 3043
rect 296686 3012 337117 3040
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 120166 2972 120172 2984
rect 116688 2944 120172 2972
rect 116581 2935 116639 2941
rect 120166 2932 120172 2944
rect 120224 2932 120230 2984
<<<<<<< HEAD
rect 291378 2932 291384 2984
rect 291436 2972 291442 2984
rect 296686 2972 296714 3012
rect 343726 3000 343732 3012
rect 343784 3000 343790 3052
=======
rect 151814 2932 151820 2984
rect 151872 2972 151878 2984
rect 160738 2972 160744 2984
rect 151872 2944 160744 2972
rect 151872 2932 151878 2944
rect 160738 2932 160744 2944
rect 160796 2932 160802 2984
rect 291378 2932 291384 2984
rect 291436 2972 291442 2984
rect 296686 2972 296714 3012
rect 337105 3009 337117 3012
rect 337151 3009 337163 3043
rect 337212 3040 337240 3080
rect 342438 3068 342444 3080
rect 342496 3068 342502 3120
rect 371142 3068 371148 3120
rect 371200 3108 371206 3120
rect 426158 3108 426164 3120
rect 371200 3080 426164 3108
rect 371200 3068 371206 3080
rect 426158 3068 426164 3080
rect 426216 3068 426222 3120
rect 431954 3068 431960 3120
rect 432012 3108 432018 3120
rect 433242 3108 433248 3120
rect 432012 3080 433248 3108
rect 432012 3068 432018 3080
rect 433242 3068 433248 3080
rect 433300 3068 433306 3120
rect 343634 3040 343640 3052
rect 337212 3012 343640 3040
rect 337105 3003 337163 3009
rect 343634 3000 343640 3012
rect 343692 3000 343698 3052
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 369762 3000 369768 3052
rect 369820 3040 369826 3052
rect 418982 3040 418988 3052
rect 369820 3012 418988 3040
rect 369820 3000 369826 3012
rect 418982 3000 418988 3012
rect 419040 3000 419046 3052
rect 291436 2944 296714 2972
rect 291436 2932 291442 2944
rect 298462 2932 298468 2984
rect 298520 2972 298526 2984
rect 299382 2972 299388 2984
rect 298520 2944 299388 2972
rect 298520 2932 298526 2944
rect 299382 2932 299388 2944
rect 299440 2932 299446 2984
rect 301958 2932 301964 2984
rect 302016 2972 302022 2984
<<<<<<< HEAD
rect 346394 2972 346400 2984
rect 302016 2944 346400 2972
rect 302016 2932 302022 2944
rect 346394 2932 346400 2944
rect 346452 2932 346458 2984
rect 351638 2932 351644 2984
rect 351696 2972 351702 2984
rect 356146 2972 356152 2984
rect 351696 2944 356152 2972
rect 351696 2932 351702 2944
rect 356146 2932 356152 2944
rect 356204 2932 356210 2984
rect 369670 2932 369676 2984
rect 369728 2972 369734 2984
rect 415486 2972 415492 2984
rect 369728 2944 415492 2972
rect 369728 2932 369734 2944
rect 415486 2932 415492 2944
rect 415544 2932 415550 2984
rect 41874 2864 41880 2916
rect 41932 2904 41938 2916
rect 42794 2904 42800 2916
rect 41932 2876 42800 2904
rect 41932 2864 41938 2876
rect 42794 2864 42800 2876
rect 42852 2864 42858 2916
=======
rect 302016 2944 345014 2972
rect 302016 2932 302022 2944
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 92750 2864 92756 2916
rect 92808 2904 92814 2916
rect 116397 2907 116455 2913
rect 116397 2904 116409 2907
rect 92808 2876 116409 2904
rect 92808 2864 92814 2876
rect 116397 2873 116409 2876
rect 116443 2873 116455 2907
rect 116397 2867 116455 2873
rect 116486 2864 116492 2916
rect 116544 2904 116550 2916
rect 119890 2904 119896 2916
rect 116544 2876 119896 2904
rect 116544 2864 116550 2876
rect 119890 2864 119896 2876
rect 119948 2864 119954 2916
rect 135438 2864 135444 2916
rect 135496 2904 135502 2916
rect 136450 2904 136456 2916
rect 135496 2876 136456 2904
rect 135496 2864 135502 2876
rect 136450 2864 136456 2876
rect 136508 2864 136514 2916
<<<<<<< HEAD
rect 190822 2864 190828 2916
rect 190880 2904 190886 2916
rect 191558 2904 191564 2916
rect 190880 2876 191564 2904
rect 190880 2864 190886 2876
rect 191558 2864 191564 2876
rect 191616 2864 191622 2916
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 220446 2864 220452 2916
rect 220504 2904 220510 2916
rect 222930 2904 222936 2916
rect 220504 2876 222936 2904
rect 220504 2864 220510 2876
rect 222930 2864 222936 2876
rect 222988 2864 222994 2916
rect 305546 2864 305552 2916
rect 305604 2904 305610 2916
<<<<<<< HEAD
rect 346486 2904 346492 2916
rect 305604 2876 346492 2904
rect 305604 2864 305610 2876
rect 346486 2864 346492 2876
rect 346544 2864 346550 2916
=======
rect 342257 2907 342315 2913
rect 342257 2904 342269 2907
rect 305604 2876 342269 2904
rect 305604 2864 305610 2876
rect 342257 2873 342269 2876
rect 342303 2873 342315 2907
rect 344986 2904 345014 2944
rect 351638 2932 351644 2984
rect 351696 2972 351702 2984
rect 356146 2972 356152 2984
rect 351696 2944 356152 2972
rect 351696 2932 351702 2944
rect 356146 2932 356152 2944
rect 356204 2932 356210 2984
rect 369670 2932 369676 2984
rect 369728 2972 369734 2984
rect 415486 2972 415492 2984
rect 369728 2944 415492 2972
rect 369728 2932 369734 2944
rect 415486 2932 415492 2944
rect 415544 2932 415550 2984
rect 346394 2904 346400 2916
rect 344986 2876 346400 2904
rect 342257 2867 342315 2873
rect 346394 2864 346400 2876
rect 346452 2864 346458 2916
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 368382 2864 368388 2916
rect 368440 2904 368446 2916
rect 368440 2876 407068 2904
rect 368440 2864 368446 2876
rect 96246 2796 96252 2848
rect 96304 2836 96310 2848
<<<<<<< HEAD
rect 96304 2808 99788 2836
rect 96304 2796 96310 2808
rect 99760 2768 99788 2808
rect 99834 2796 99840 2848
rect 99892 2836 99898 2848
rect 100294 2836 100300 2848
rect 99892 2808 100300 2836
rect 99892 2796 99898 2808
rect 100294 2796 100300 2808
rect 100352 2796 100358 2848
rect 122926 2836 122932 2848
rect 100404 2808 122932 2836
rect 100404 2768 100432 2808
=======
rect 122926 2836 122932 2848
rect 96304 2808 122932 2836
rect 96304 2796 96310 2808
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 122926 2796 122932 2808
rect 122984 2796 122990 2848
rect 309042 2796 309048 2848
rect 309100 2836 309106 2848
rect 347958 2836 347964 2848
rect 309100 2808 347964 2836
rect 309100 2796 309106 2808
rect 347958 2796 347964 2808
rect 348016 2796 348022 2848
rect 366910 2796 366916 2848
rect 366968 2836 366974 2848
rect 404814 2836 404820 2848
rect 366968 2808 404820 2836
rect 366968 2796 366974 2808
rect 404814 2796 404820 2808
rect 404872 2796 404878 2848
rect 407040 2836 407068 2876
rect 407114 2864 407120 2916
rect 407172 2904 407178 2916
rect 408402 2904 408408 2916
rect 407172 2876 408408 2904
rect 407172 2864 407178 2876
rect 408402 2864 408408 2876
rect 408460 2864 408466 2916
rect 411898 2836 411904 2848
rect 407040 2808 411904 2836
rect 411898 2796 411904 2808
rect 411956 2796 411962 2848
<<<<<<< HEAD
rect 99760 2740 100432 2768
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
<< via1 >>
rect 315948 700952 316000 701004
rect 413652 700952 413704 701004
rect 325608 700884 325660 700936
rect 429844 700884 429896 700936
rect 335268 700816 335320 700868
rect 446128 700816 446180 700868
rect 346308 700748 346360 700800
rect 462320 700748 462372 700800
rect 256608 700680 256660 700732
rect 316316 700680 316368 700732
rect 355968 700680 356020 700732
rect 478512 700680 478564 700732
rect 267556 700612 267608 700664
rect 332508 700612 332560 700664
rect 365628 700612 365680 700664
rect 494796 700612 494848 700664
rect 217968 700544 218020 700596
rect 251456 700544 251508 700596
rect 277308 700544 277360 700596
rect 348792 700544 348844 700596
rect 375288 700544 375340 700596
rect 510988 700544 511040 700596
rect 227628 700476 227680 700528
rect 267648 700476 267700 700528
rect 286968 700476 287020 700528
rect 364984 700476 365036 700528
rect 384948 700476 385000 700528
rect 527180 700476 527232 700528
rect 188988 700408 189040 700460
rect 202788 700408 202840 700460
rect 237288 700408 237340 700460
rect 283840 700408 283892 700460
rect 296628 700408 296680 700460
rect 381176 700408 381228 700460
rect 394608 700408 394660 700460
rect 543464 700408 543516 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 56784 700340 56836 700392
rect 71044 700340 71096 700392
rect 177948 700340 178000 700392
rect 186504 700340 186556 700392
rect 198648 700340 198700 700392
rect 218980 700340 219032 700392
rect 220084 700340 220136 700392
rect 235172 700340 235224 700392
rect 246948 700340 247000 700392
rect 300124 700340 300176 700392
rect 306288 700340 306340 700392
rect 397460 700340 397512 700392
rect 404268 700340 404320 700392
rect 559656 700340 559708 700392
rect 62028 700272 62080 700324
rect 575848 700272 575900 700324
rect 121644 700204 121696 700256
rect 122748 700204 122800 700256
rect 154120 700068 154172 700120
rect 155224 700068 155276 700120
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 169024 699660 169076 699712
rect 170312 699660 170364 699712
rect 411904 696940 411956 696992
rect 580172 696940 580224 696992
rect 3148 683136 3200 683188
rect 11704 683136 11756 683188
rect 406384 683136 406436 683188
rect 580172 683136 580224 683188
rect 406476 670692 406528 670744
rect 580172 670692 580224 670744
rect 3148 656888 3200 656940
rect 22744 656888 22796 656940
rect 410524 643084 410576 643136
rect 580172 643084 580224 643136
rect 3332 632068 3384 632120
rect 14464 632068 14516 632120
rect 418804 630640 418856 630692
rect 579988 630640 580040 630692
rect 2964 618264 3016 618316
rect 35164 618264 35216 618316
rect 406568 616836 406620 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 25504 605820 25556 605872
rect 2780 592288 2832 592340
rect 4804 592288 4856 592340
rect 406660 590656 406712 590708
rect 579620 590656 579672 590708
rect 3332 579640 3384 579692
rect 15844 579640 15896 579692
rect 406752 576852 406804 576904
rect 579620 576852 579672 576904
rect 3056 565836 3108 565888
rect 36544 565836 36596 565888
rect 406844 563048 406896 563100
rect 579896 563048 579948 563100
rect 3332 553392 3384 553444
rect 29644 553392 29696 553444
rect 3332 539656 3384 539708
rect 7564 539656 7616 539708
rect 407764 536800 407816 536852
rect 580172 536800 580224 536852
rect 3332 527144 3384 527196
rect 17224 527144 17276 527196
rect 417424 524424 417476 524476
rect 580172 524424 580224 524476
rect 3240 500964 3292 501016
rect 32404 500964 32456 501016
rect 406936 484372 406988 484424
rect 579620 484372 579672 484424
rect 2872 474716 2924 474768
rect 18604 474716 18656 474768
rect 407028 470568 407080 470620
rect 579988 470568 580040 470620
rect 3056 462340 3108 462392
rect 39304 462340 39356 462392
rect 2964 448536 3016 448588
rect 33784 448536 33836 448588
rect 414664 430584 414716 430636
rect 579988 430584 580040 430636
rect 2964 422288 3016 422340
rect 21364 422288 21416 422340
rect 406292 418140 406344 418192
rect 580172 418140 580224 418192
rect 406200 404336 406252 404388
rect 580172 404336 580224 404388
rect 406108 378156 406160 378208
rect 579804 378156 579856 378208
rect 60832 369792 60884 369844
rect 62028 369792 62080 369844
rect 168104 369792 168156 369844
rect 169024 369792 169076 369844
rect 217232 369792 217284 369844
rect 217968 369792 218020 369844
rect 227076 369792 227128 369844
rect 227628 369792 227680 369844
rect 286048 369792 286100 369844
rect 286968 369792 287020 369844
rect 295892 369792 295944 369844
rect 296628 369792 296680 369844
rect 305736 369792 305788 369844
rect 306288 369792 306340 369844
rect 354864 369792 354916 369844
rect 355968 369792 356020 369844
rect 364708 369792 364760 369844
rect 365628 369792 365680 369844
rect 374552 369792 374604 369844
rect 375288 369792 375340 369844
rect 384396 369792 384448 369844
rect 384948 369792 385000 369844
rect 402980 369792 403032 369844
rect 404268 369792 404320 369844
rect 197636 369656 197688 369708
rect 198648 369656 198700 369708
rect 71044 369316 71096 369368
rect 99288 369316 99340 369368
rect 41328 369248 41380 369300
rect 89444 369248 89496 369300
rect 106188 369248 106240 369300
rect 128820 369248 128872 369300
rect 24768 369180 24820 369232
rect 79600 369180 79652 369232
rect 89628 369180 89680 369232
rect 118976 369180 119028 369232
rect 137928 369180 137980 369232
rect 148416 369180 148468 369232
rect 155224 369180 155276 369232
rect 158260 369180 158312 369232
rect 8208 369112 8260 369164
rect 69756 369112 69808 369164
rect 73068 369112 73120 369164
rect 109132 369112 109184 369164
rect 122748 369112 122800 369164
rect 138572 369112 138624 369164
rect 187792 369112 187844 369164
rect 188988 369112 189040 369164
rect 207480 369112 207532 369164
rect 220084 369112 220136 369164
rect 345112 369112 345164 369164
rect 346308 369112 346360 369164
rect 266452 369044 266504 369096
rect 267648 369044 267700 369096
rect 276296 368976 276348 369028
rect 277308 368976 277360 369028
rect 3424 365644 3476 365696
rect 57428 365644 57480 365696
rect 406016 364964 406068 365016
rect 411904 364964 411956 365016
rect 411996 364352 412048 364404
rect 580172 364352 580224 364404
rect 11704 361496 11756 361548
rect 57152 361496 57204 361548
rect 3516 355988 3568 356040
rect 57244 355988 57296 356040
rect 406384 351908 406436 351960
rect 580172 351908 580224 351960
rect 22744 350480 22796 350532
rect 57612 350480 57664 350532
rect 406476 349052 406528 349104
rect 580080 349052 580132 349104
rect 3608 344972 3660 345024
rect 57612 344972 57664 345024
rect 406476 343340 406528 343392
rect 410524 343340 410576 343392
rect 14464 339396 14516 339448
rect 57612 339396 57664 339448
rect 406476 338036 406528 338088
rect 418804 338036 418856 338088
rect 35164 333888 35216 333940
rect 57612 333888 57664 333940
rect 25504 328380 25556 328432
rect 57336 328380 57388 328432
rect 406568 327020 406620 327072
rect 580356 327020 580408 327072
rect 406476 324300 406528 324352
rect 580172 324300 580224 324352
rect 4804 322872 4856 322924
rect 57336 322872 57388 322924
rect 15844 317364 15896 317416
rect 57612 317364 57664 317416
rect 406568 311856 406620 311908
rect 580172 311856 580224 311908
rect 36544 310428 36596 310480
rect 57612 310428 57664 310480
rect 29644 304920 29696 304972
rect 57428 304920 57480 304972
rect 406844 304920 406896 304972
rect 580448 304920 580500 304972
rect 7564 299412 7616 299464
rect 57612 299412 57664 299464
rect 405832 299276 405884 299328
rect 407764 299276 407816 299328
rect 406660 298120 406712 298172
rect 580172 298120 580224 298172
rect 17224 293904 17276 293956
rect 57612 293904 57664 293956
rect 406844 292476 406896 292528
rect 417424 292476 417476 292528
rect 3700 288328 3752 288380
rect 57612 288328 57664 288380
rect 406844 286968 406896 287020
rect 580540 286968 580592 287020
rect 32404 282820 32456 282872
rect 57612 282820 57664 282872
rect 406844 281460 406896 281512
rect 580632 281460 580684 281512
rect 3792 277312 3844 277364
rect 57612 277312 57664 277364
rect 406752 271872 406804 271924
rect 580172 271872 580224 271924
rect 18604 271804 18656 271856
rect 57520 271804 57572 271856
rect 39304 266296 39356 266348
rect 57336 266296 57388 266348
rect 407028 264868 407080 264920
rect 580724 264868 580776 264920
rect 33784 260788 33836 260840
rect 57428 260788 57480 260840
rect 406936 259360 406988 259412
rect 580816 259360 580868 259412
rect 406844 258068 406896 258120
rect 580172 258068 580224 258120
rect 3884 255212 3936 255264
rect 57612 255212 57664 255264
rect 407028 252832 407080 252884
rect 414664 252832 414716 252884
rect 21364 249704 21416 249756
rect 57244 249704 57296 249756
rect 406936 244264 406988 244316
rect 580172 244264 580224 244316
rect 3976 244196 4028 244248
rect 57428 244196 57480 244248
rect 4068 238688 4120 238740
rect 57612 238688 57664 238740
rect 407028 235900 407080 235952
rect 580908 235900 580960 235952
rect 3332 233180 3384 233232
rect 57612 233180 57664 233232
rect 407028 231820 407080 231872
rect 579620 231820 579672 231872
rect 3240 227672 3292 227724
rect 57612 227672 57664 227724
rect 406292 224612 406344 224664
rect 411996 224612 412048 224664
rect 3424 222096 3476 222148
rect 57612 222096 57664 222148
rect 406292 218016 406344 218068
rect 580172 218016 580224 218068
rect 3516 216588 3568 216640
rect 57060 216588 57112 216640
rect 406384 213868 406436 213920
rect 580264 213868 580316 213920
rect 3608 211080 3660 211132
rect 56784 211080 56836 211132
rect 406384 205640 406436 205692
rect 580172 205640 580224 205692
rect 3148 205572 3200 205624
rect 57612 205572 57664 205624
rect 3056 200064 3108 200116
rect 57612 200064 57664 200116
rect 2964 194488 3016 194540
rect 57612 194488 57664 194540
rect 406476 191836 406528 191888
rect 580172 191836 580224 191888
rect 406752 191768 406804 191820
rect 580356 191768 580408 191820
rect 3700 188980 3752 189032
rect 57612 188980 57664 189032
rect 3792 183472 3844 183524
rect 57612 183472 57664 183524
rect 406568 178032 406620 178084
rect 580172 178032 580224 178084
rect 2872 177964 2924 178016
rect 56692 177964 56744 178016
rect 3884 172456 3936 172508
rect 57612 172456 57664 172508
rect 3976 166948 4028 167000
rect 57612 166948 57664 167000
rect 406660 165588 406712 165640
rect 580172 165588 580224 165640
rect 3424 161372 3476 161424
rect 57612 161372 57664 161424
rect 3516 155864 3568 155916
rect 57612 155864 57664 155916
rect 406384 151784 406436 151836
rect 579988 151784 580040 151836
rect 3608 150356 3660 150408
rect 56876 150356 56928 150408
rect 3700 144848 3752 144900
rect 57520 144848 57572 144900
rect 3792 139340 3844 139392
rect 57520 139340 57572 139392
rect 406476 137980 406528 138032
rect 580172 137980 580224 138032
rect 3424 133832 3476 133884
rect 57520 133832 57572 133884
rect 3516 128256 3568 128308
rect 56968 128256 57020 128308
rect 407028 125604 407080 125656
rect 580172 125604 580224 125656
rect 3608 122748 3660 122800
rect 57060 122748 57112 122800
rect 3424 115948 3476 116000
rect 57612 115948 57664 116000
rect 406384 113092 406436 113144
rect 579804 113092 579856 113144
rect 3516 110440 3568 110492
rect 57612 110440 57664 110492
rect 3424 104864 3476 104916
rect 57428 104864 57480 104916
rect 406476 100648 406528 100700
rect 580172 100648 580224 100700
rect 3884 99356 3936 99408
rect 57428 99356 57480 99408
rect 3792 93848 3844 93900
rect 57612 93848 57664 93900
rect 3700 88340 3752 88392
rect 57520 88340 57572 88392
rect 406384 86912 406436 86964
rect 580172 86912 580224 86964
rect 3608 82832 3660 82884
rect 57428 82832 57480 82884
rect 3516 77256 3568 77308
rect 57520 77256 57572 77308
rect 406844 73108 406896 73160
rect 580172 73108 580224 73160
rect 3424 71748 3476 71800
rect 57428 71748 57480 71800
rect 60832 71748 60884 71800
rect 62067 71748 62119 71800
rect 98000 71748 98052 71800
rect 99051 71748 99103 71800
rect 100760 71748 100812 71800
rect 101842 71748 101894 71800
rect 109132 71748 109184 71800
rect 110216 71748 110268 71800
rect 114560 71748 114612 71800
rect 115798 71748 115850 71800
rect 116032 71748 116084 71800
rect 117194 71748 117246 71800
rect 117320 71748 117372 71800
rect 118589 71748 118641 71800
rect 118792 71748 118844 71800
rect 119985 71748 120037 71800
rect 120172 71748 120224 71800
rect 121380 71748 121432 71800
rect 230480 71748 230532 71800
rect 231633 71748 231685 71800
rect 234712 71748 234764 71800
rect 235820 71748 235872 71800
rect 236092 71748 236144 71800
rect 237215 71748 237267 71800
rect 237380 71748 237432 71800
rect 238611 71748 238663 71800
rect 240140 71748 240192 71800
rect 241402 71748 241454 71800
rect 321560 71748 321612 71800
rect 322347 71748 322399 71800
rect 324320 71748 324372 71800
rect 325138 71748 325190 71800
rect 327080 71748 327132 71800
rect 327929 71748 327981 71800
rect 328460 71748 328512 71800
rect 329325 71748 329377 71800
rect 329840 71748 329892 71800
rect 330720 71748 330772 71800
rect 331220 71748 331272 71800
rect 332116 71748 332168 71800
rect 333980 71748 334032 71800
rect 334907 71748 334959 71800
rect 335452 71748 335504 71800
rect 336303 71748 336355 71800
rect 338120 71748 338172 71800
rect 339094 71748 339146 71800
rect 340972 71748 341024 71800
rect 341885 71748 341937 71800
rect 349252 71748 349304 71800
rect 350259 71748 350311 71800
rect 53104 70320 53156 70372
rect 64144 70320 64196 70372
rect 148968 70320 149020 70372
rect 227444 70320 227496 70372
rect 265808 70320 265860 70372
<<<<<<< HEAD
rect 295984 70320 296036 70372
rect 299388 70320 299440 70372
rect 346032 70320 346084 70372
rect 375380 70320 375432 70372
rect 447140 70320 447192 70372
=======
rect 295892 70320 295944 70372
rect 299388 70320 299440 70372
rect 346032 70320 346084 70372
rect 374000 70320 374052 70372
rect 440240 70320 440292 70372
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 41328 70252 41380 70304
rect 67640 70252 67692 70304
rect 121368 70252 121420 70304
rect 128360 70252 128412 70304
rect 141976 70252 142028 70304
rect 226064 70252 226116 70304
<<<<<<< HEAD
rect 287704 70252 287756 70304
rect 325792 70252 325844 70304
rect 338028 70252 338080 70304
rect 353760 70252 353812 70304
rect 378232 70252 378284 70304
=======
rect 294420 70252 294472 70304
rect 295984 70252 296036 70304
rect 325792 70252 325844 70304
rect 338028 70252 338080 70304
rect 353760 70252 353812 70304
rect 375380 70252 375432 70304
rect 447140 70252 447192 70304
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 34428 70184 34480 70236
rect 64880 70184 64932 70236
rect 50344 70116 50396 70168
rect 84384 70184 84436 70236
rect 119344 70184 119396 70236
rect 127624 70184 127676 70236
rect 144828 70184 144880 70236
rect 226708 70184 226760 70236
rect 291660 70184 291712 70236
rect 345388 70184 345440 70236
<<<<<<< HEAD
rect 380992 70184 381044 70236
rect 454040 70252 454092 70304
rect 460940 70184 460992 70236
=======
rect 379612 70184 379664 70236
rect 454040 70184 454092 70236
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 80888 70116 80940 70168
rect 27528 70048 27580 70100
rect 68284 70048 68336 70100
rect 95516 70116 95568 70168
rect 106740 70116 106792 70168
rect 122840 70116 122892 70168
rect 137928 70116 137980 70168
rect 225328 70116 225380 70168
rect 231124 70116 231176 70168
rect 239956 70116 240008 70168
<<<<<<< HEAD
rect 281448 70116 281500 70168
rect 342352 70116 342404 70168
rect 379612 70116 379664 70168
rect 467840 70116 467892 70168
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 103428 70048 103480 70100
rect 107476 70048 107528 70100
rect 125600 70048 125652 70100
rect 163964 70048 164016 70100
<<<<<<< HEAD
rect 250352 70048 250404 70100
=======
rect 250352 70116 250404 70168
rect 281448 70116 281500 70168
rect 342352 70116 342404 70168
rect 378232 70116 378284 70168
rect 460940 70116 460992 70168
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 295800 70048 295852 70100
rect 410524 70048 410576 70100
rect 51724 69980 51776 70032
rect 92020 69980 92072 70032
rect 124864 69980 124916 70032
rect 135168 69980 135220 70032
rect 224684 69980 224736 70032
rect 234528 69980 234580 70032
rect 244188 69980 244240 70032
rect 295156 69980 295208 70032
rect 418804 69980 418856 70032
rect 17868 69912 17920 69964
rect 63500 69912 63552 69964
rect 107568 69912 107620 69964
rect 114468 69912 114520 69964
rect 126980 69912 127032 69964
rect 353944 69912 353996 69964
<<<<<<< HEAD
rect 474740 69912 474792 69964
=======
rect 380992 69912 381044 69964
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 7564 69844 7616 69896
rect 60280 69844 60332 69896
rect 65524 69844 65576 69896
rect 92480 69844 92532 69896
rect 93124 69844 93176 69896
rect 94136 69844 94188 69896
rect 103244 69844 103296 69896
rect 104164 69844 104216 69896
rect 124128 69844 124180 69896
<<<<<<< HEAD
rect 131028 69844 131080 69896
rect 223948 69844 224000 69896
rect 228364 69844 228416 69896
rect 230204 69844 230256 69896
rect 242808 69844 242860 69896
rect 250444 69844 250496 69896
rect 264980 69844 265032 69896
rect 472624 69844 472676 69896
=======
rect 129648 69844 129700 69896
rect 134616 69844 134668 69896
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 18604 69776 18656 69828
rect 107660 69776 107712 69828
rect 111708 69776 111760 69828
rect 126244 69776 126296 69828
<<<<<<< HEAD
rect 129648 69776 129700 69828
rect 134616 69776 134668 69828
rect 154212 69776 154264 69828
rect 204996 69776 205048 69828
rect 208584 69776 208636 69828
rect 413284 69776 413336 69828
rect 21364 69708 21416 69760
rect 130476 69708 130528 69760
rect 411904 69708 411956 69760
=======
rect 131028 69776 131080 69828
rect 371792 69844 371844 69896
rect 467840 69912 467892 69964
rect 474740 69844 474792 69896
rect 223948 69776 224000 69828
rect 228364 69776 228416 69828
rect 230204 69776 230256 69828
rect 242808 69776 242860 69828
rect 250444 69776 250496 69828
rect 264980 69776 265032 69828
rect 287704 69776 287756 69828
rect 472624 69776 472676 69828
rect 21364 69708 21416 69760
rect 130476 69708 130528 69760
rect 154212 69708 154264 69760
rect 204904 69708 204956 69760
rect 208584 69708 208636 69760
rect 413284 69708 413336 69760
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 11704 69640 11756 69692
rect 133236 69640 133288 69692
rect 193312 69640 193364 69692
rect 205088 69640 205140 69692
<<<<<<< HEAD
rect 371792 69640 371844 69692
rect 376760 69640 376812 69692
=======
rect 411904 69640 411956 69692
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 66260 69572 66312 69624
rect 81624 69572 81676 69624
rect 86224 69572 86276 69624
rect 100668 69572 100720 69624
rect 155868 69572 155920 69624
rect 65892 69504 65944 69556
rect 66904 69504 66956 69556
rect 157708 69504 157760 69556
rect 224224 69504 224276 69556
rect 227628 69572 227680 69624
rect 247684 69572 247736 69624
rect 248972 69572 249024 69624
<<<<<<< HEAD
rect 272156 69572 272208 69624
rect 274364 69572 274416 69624
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 293776 69572 293828 69624
rect 310152 69572 310204 69624
rect 313188 69572 313240 69624
rect 348884 69572 348936 69624
<<<<<<< HEAD
rect 374000 69572 374052 69624
rect 440240 69572 440292 69624
=======
rect 372620 69572 372672 69624
rect 431960 69572 432012 69624
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 228824 69504 228876 69556
rect 291844 69504 291896 69556
rect 323032 69504 323084 69556
rect 324228 69504 324280 69556
rect 350632 69504 350684 69556
<<<<<<< HEAD
rect 372620 69504 372672 69556
rect 431960 69504 432012 69556
rect 164700 69436 164752 69488
rect 226984 69436 227036 69488
=======
rect 371884 69504 371936 69556
rect 429200 69504 429252 69556
rect 164700 69436 164752 69488
rect 226984 69436 227036 69488
rect 272156 69436 272208 69488
rect 274364 69436 274416 69488
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 289084 69436 289136 69488
rect 320272 69436 320324 69488
rect 342168 69436 342220 69488
rect 354404 69436 354456 69488
<<<<<<< HEAD
rect 371884 69436 371936 69488
rect 429200 69436 429252 69488
=======
rect 370504 69436 370556 69488
rect 422300 69436 422352 69488
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 126888 69368 126940 69420
rect 133880 69368 133932 69420
rect 154856 69368 154908 69420
rect 206284 69368 206336 69420
rect 209688 69368 209740 69420
rect 239312 69368 239364 69420
rect 293040 69368 293092 69420
rect 310336 69368 310388 69420
<<<<<<< HEAD
rect 370504 69368 370556 69420
rect 422300 69368 422352 69420
=======
rect 367744 69368 367796 69420
rect 407120 69368 407172 69420
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 156328 69300 156380 69352
rect 204904 69300 204956 69352
rect 207204 69300 207256 69352
rect 224316 69300 224368 69352
rect 290280 69300 290332 69352
rect 292396 69300 292448 69352
rect 295248 69300 295300 69352
<<<<<<< HEAD
rect 367744 69300 367796 69352
rect 407120 69300 407172 69352
=======
rect 376760 69300 376812 69352
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 111800 69232 111852 69284
rect 114376 69232 114428 69284
rect 163228 69232 163280 69284
rect 209136 69232 209188 69284
rect 222844 69232 222896 69284
rect 233240 69232 233292 69284
<<<<<<< HEAD
rect 294420 69232 294472 69284
rect 295892 69232 295944 69284
rect 309876 69232 309928 69284
rect 319536 69232 319588 69284
rect 383752 69232 383804 69284
rect 414664 69232 414716 69284
=======
rect 309876 69232 309928 69284
rect 319536 69232 319588 69284
rect 383752 69232 383804 69284
rect 414664 69300 414716 69352
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 78128 69164 78180 69216
rect 83464 69164 83516 69216
rect 198004 69164 198056 69216
rect 236460 69164 236512 69216
rect 57244 69096 57296 69148
rect 61384 69096 61436 69148
rect 72424 69096 72476 69148
rect 73252 69096 73304 69148
rect 74632 69096 74684 69148
rect 75736 69096 75788 69148
rect 76012 69096 76064 69148
rect 77116 69096 77168 69148
rect 78864 69096 78916 69148
rect 79968 69096 80020 69148
rect 94504 69096 94556 69148
rect 100392 69096 100444 69148
rect 173072 69096 173124 69148
rect 173808 69096 173860 69148
rect 186320 69096 186372 69148
rect 187608 69096 187660 69148
rect 187700 69096 187752 69148
rect 188896 69096 188948 69148
rect 189080 69096 189132 69148
rect 190276 69096 190328 69148
rect 190460 69096 190512 69148
rect 191656 69096 191708 69148
rect 194692 69096 194744 69148
rect 195888 69096 195940 69148
rect 196072 69096 196124 69148
rect 197176 69096 197228 69148
rect 198832 69096 198884 69148
rect 199936 69096 199988 69148
rect 203708 69096 203760 69148
rect 58624 69028 58676 69080
rect 60648 69028 60700 69080
rect 69664 69028 69716 69080
rect 71780 69028 71832 69080
rect 73068 69028 73120 69080
rect 73896 69028 73948 69080
rect 75368 69028 75420 69080
rect 75828 69028 75880 69080
rect 76748 69028 76800 69080
rect 77208 69028 77260 69080
rect 77392 69028 77444 69080
rect 79324 69028 79376 69080
rect 80244 69028 80296 69080
rect 81348 69028 81400 69080
rect 83004 69028 83056 69080
rect 84108 69028 84160 69080
rect 87604 69028 87656 69080
rect 91376 69028 91428 69080
rect 94596 69028 94648 69080
rect 96252 69028 96304 69080
rect 98644 69028 98696 69080
rect 99748 69028 99800 69080
rect 103980 69028 104032 69080
rect 104808 69028 104860 69080
rect 105360 69028 105412 69080
rect 106096 69028 106148 69080
rect 125508 69028 125560 69080
rect 129004 69028 129056 69080
rect 133788 69028 133840 69080
rect 135352 69028 135404 69080
rect 136732 69028 136784 69080
rect 137836 69028 137888 69080
rect 138112 69028 138164 69080
rect 139308 69028 139360 69080
rect 139584 69028 139636 69080
rect 140688 69028 140740 69080
rect 140964 69028 141016 69080
rect 142068 69028 142120 69080
rect 142344 69028 142396 69080
rect 143448 69028 143500 69080
rect 143724 69028 143776 69080
rect 144644 69028 144696 69080
rect 145104 69028 145156 69080
rect 146116 69028 146168 69080
rect 146484 69028 146536 69080
rect 147588 69028 147640 69080
rect 147956 69028 148008 69080
rect 148876 69028 148928 69080
rect 149336 69028 149388 69080
rect 150256 69028 150308 69080
rect 150716 69028 150768 69080
rect 151728 69028 151780 69080
rect 152096 69028 152148 69080
rect 153016 69028 153068 69080
rect 153476 69028 153528 69080
rect 154488 69028 154540 69080
rect 159088 69028 159140 69080
rect 159916 69028 159968 69080
rect 160468 69028 160520 69080
rect 161388 69028 161440 69080
rect 161848 69028 161900 69080
rect 162676 69028 162728 69080
rect 166080 69028 166132 69080
rect 166816 69028 166868 69080
rect 167460 69028 167512 69080
rect 168288 69028 168340 69080
rect 168840 69028 168892 69080
rect 169668 69028 169720 69080
rect 170220 69028 170272 69080
rect 170956 69028 171008 69080
rect 171600 69028 171652 69080
rect 173164 69028 173216 69080
rect 174452 69028 174504 69080
rect 175096 69028 175148 69080
rect 175832 69028 175884 69080
rect 176476 69028 176528 69080
rect 178592 69028 178644 69080
rect 179236 69028 179288 69080
rect 179972 69028 180024 69080
rect 180616 69028 180668 69080
rect 181444 69028 181496 69080
rect 182088 69028 182140 69080
rect 182824 69028 182876 69080
rect 183376 69028 183428 69080
rect 184204 69028 184256 69080
rect 184848 69028 184900 69080
rect 185584 69028 185636 69080
rect 186228 69028 186280 69080
rect 186964 69028 187016 69080
rect 187516 69028 187568 69080
rect 188344 69028 188396 69080
rect 188988 69028 189040 69080
rect 189816 69028 189868 69080
rect 190368 69028 190420 69080
rect 191196 69028 191248 69080
rect 191748 69028 191800 69080
rect 191840 69028 191892 69080
rect 193128 69028 193180 69080
rect 195336 69028 195388 69080
rect 195796 69028 195848 69080
rect 196716 69028 196768 69080
rect 197268 69028 197320 69080
rect 198188 69028 198240 69080
rect 198648 69028 198700 69080
rect 199568 69028 199620 69080
rect 200028 69028 200080 69080
rect 200212 69028 200264 69080
rect 201408 69028 201460 69080
rect 201684 69028 201736 69080
rect 202788 69028 202840 69080
rect 203064 69028 203116 69080
rect 204168 69028 204220 69080
rect 207940 69096 207992 69148
<<<<<<< HEAD
rect 213552 69096 213604 69148
=======
rect 213644 69096 213696 69148
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 248420 69096 248472 69148
rect 249708 69096 249760 69148
rect 251180 69096 251232 69148
rect 252468 69096 252520 69148
rect 252560 69096 252612 69148
rect 253848 69096 253900 69148
rect 253940 69096 253992 69148
rect 255228 69096 255280 69148
rect 255412 69096 255464 69148
rect 256608 69096 256660 69148
rect 256792 69096 256844 69148
rect 257896 69096 257948 69148
rect 258172 69096 258224 69148
rect 259276 69096 259328 69148
rect 260932 69096 260984 69148
rect 262036 69096 262088 69148
rect 262312 69096 262364 69148
rect 263416 69096 263468 69148
rect 310520 69096 310572 69148
rect 311808 69096 311860 69148
rect 327724 69096 327776 69148
rect 332784 69096 332836 69148
rect 389364 69096 389416 69148
rect 390376 69096 390428 69148
<<<<<<< HEAD
rect 390744 69096 390796 69148
rect 392400 69096 392452 69148
rect 403348 69096 403400 69148
rect 404176 69096 404228 69148
=======
rect 401876 69096 401928 69148
rect 403716 69096 403768 69148
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 210056 69028 210108 69080
rect 210976 69028 211028 69080
rect 211436 69028 211488 69080
rect 212356 69028 212408 69080
rect 212816 69028 212868 69080
rect 213828 69028 213880 69080
rect 214196 69028 214248 69080
rect 215116 69028 215168 69080
rect 215576 69028 215628 69080
rect 216496 69028 216548 69080
rect 216956 69028 217008 69080
rect 217876 69028 217928 69080
rect 218428 69028 218480 69080
rect 218980 69028 219032 69080
rect 219808 69028 219860 69080
rect 220636 69028 220688 69080
rect 221188 69028 221240 69080
rect 222108 69028 222160 69080
rect 232504 69028 232556 69080
rect 235080 69028 235132 69080
rect 242164 69028 242216 69080
rect 243452 69028 243504 69080
rect 249064 69028 249116 69080
rect 249616 69028 249668 69080
rect 249800 69028 249852 69080
rect 251088 69028 251140 69080
rect 251916 69028 251968 69080
rect 252376 69028 252428 69080
rect 253296 69028 253348 69080
rect 253756 69028 253808 69080
rect 254676 69028 254728 69080
rect 255136 69028 255188 69080
rect 256056 69028 256108 69080
rect 256516 69028 256568 69080
rect 257436 69028 257488 69080
rect 257988 69028 258040 69080
rect 258908 69028 258960 69080
rect 259368 69028 259420 69080
rect 259552 69028 259604 69080
rect 260748 69028 260800 69080
rect 261668 69028 261720 69080
rect 262128 69028 262180 69080
rect 263048 69028 263100 69080
rect 263508 69028 263560 69080
rect 263784 69028 263836 69080
rect 264888 69028 264940 69080
rect 265164 69028 265216 69080
rect 266268 69028 266320 69080
rect 266544 69028 266596 69080
rect 267648 69028 267700 69080
rect 267924 69028 267976 69080
rect 269028 69028 269080 69080
rect 269304 69028 269356 69080
rect 270316 69028 270368 69080
rect 270684 69028 270736 69080
rect 271696 69028 271748 69080
rect 273536 69028 273588 69080
rect 274456 69028 274508 69080
rect 274916 69028 274968 69080
rect 275836 69028 275888 69080
rect 276296 69028 276348 69080
rect 277216 69028 277268 69080
rect 277676 69028 277728 69080
rect 278596 69028 278648 69080
rect 279056 69028 279108 69080
rect 279976 69028 280028 69080
rect 280528 69028 280580 69080
rect 281356 69028 281408 69080
rect 281908 69028 281960 69080
rect 282736 69028 282788 69080
rect 283288 69028 283340 69080
rect 284208 69028 284260 69080
rect 284668 69028 284720 69080
rect 285496 69028 285548 69080
rect 286048 69028 286100 69080
rect 286876 69028 286928 69080
rect 287428 69028 287480 69080
rect 288348 69028 288400 69080
rect 288900 69028 288952 69080
rect 289728 69028 289780 69080
rect 290924 69028 290976 69080
rect 293776 69028 293828 69080
rect 297272 69028 297324 69080
rect 298008 69028 298060 69080
rect 298652 69028 298704 69080
rect 299296 69028 299348 69080
rect 300032 69028 300084 69080
rect 300676 69028 300728 69080
rect 301412 69028 301464 69080
rect 302148 69028 302200 69080
rect 302792 69028 302844 69080
rect 303528 69028 303580 69080
rect 304264 69028 304316 69080
rect 304816 69028 304868 69080
rect 305644 69028 305696 69080
rect 306196 69028 306248 69080
rect 307024 69028 307076 69080
rect 307668 69028 307720 69080
rect 308404 69028 308456 69080
rect 309048 69028 309100 69080
rect 309784 69028 309836 69080
rect 310428 69028 310480 69080
rect 311164 69028 311216 69080
rect 311716 69028 311768 69080
rect 311900 69028 311952 69080
rect 313096 69028 313148 69080
rect 331864 69028 331916 69080
rect 333520 69028 333572 69080
rect 359372 69028 359424 69080
rect 360108 69028 360160 69080
rect 360752 69028 360804 69080
rect 361396 69028 361448 69080
rect 362132 69028 362184 69080
rect 362868 69028 362920 69080
rect 363512 69028 363564 69080
rect 364248 69028 364300 69080
rect 364892 69028 364944 69080
rect 365628 69028 365680 69080
rect 366364 69028 366416 69080
rect 366916 69028 366968 69080
rect 369124 69028 369176 69080
rect 369676 69028 369728 69080
rect 373264 69028 373316 69080
rect 373908 69028 373960 69080
rect 374736 69028 374788 69080
rect 375288 69028 375340 69080
rect 376116 69028 376168 69080
rect 376668 69028 376720 69080
rect 377496 69028 377548 69080
rect 378048 69028 378100 69080
rect 378876 69028 378928 69080
rect 379428 69028 379480 69080
rect 380256 69028 380308 69080
rect 380808 69028 380860 69080
rect 381636 69028 381688 69080
rect 382188 69028 382240 69080
rect 382372 69028 382424 69080
rect 383568 69028 383620 69080
rect 385868 69028 385920 69080
rect 386328 69028 386380 69080
rect 388628 69028 388680 69080
rect 389088 69028 389140 69080
rect 390008 69028 390060 69080
rect 390468 69028 390520 69080
<<<<<<< HEAD
=======
rect 390744 69028 390796 69080
rect 391940 69028 391992 69080
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 392124 69028 392176 69080
rect 393136 69028 393188 69080
rect 393504 69028 393556 69080
rect 394516 69028 394568 69080
rect 394976 69028 395028 69080
rect 395896 69028 395948 69080
rect 396356 69028 396408 69080
rect 397276 69028 397328 69080
rect 397736 69028 397788 69080
rect 398748 69028 398800 69080
rect 399116 69028 399168 69080
rect 400128 69028 400180 69080
rect 400496 69028 400548 69080
rect 401508 69028 401560 69080
<<<<<<< HEAD
rect 401876 69028 401928 69080
=======
rect 403348 69028 403400 69080
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 404268 69028 404320 69080
rect 384488 68824 384540 68876
rect 492680 68824 492732 68876
rect 55128 68756 55180 68808
rect 70400 68756 70452 68808
rect 172336 68756 172388 68808
rect 320180 68756 320232 68808
rect 386604 68756 386656 68808
rect 503720 68756 503772 68808
rect 48228 68688 48280 68740
rect 69020 68688 69072 68740
rect 177212 68688 177264 68740
rect 345020 68688 345072 68740
rect 391480 68688 391532 68740
rect 528560 68688 528612 68740
rect 37188 68620 37240 68672
rect 65892 68620 65944 68672
rect 310336 68620 310388 68672
rect 481640 68620 481692 68672
rect 14464 68552 14516 68604
rect 62764 68552 62816 68604
<<<<<<< HEAD
rect 177304 68552 177356 68604
rect 229560 68552 229612 68604
rect 244372 68552 244424 68604
rect 245568 68552 245620 68604
rect 295892 68552 295944 68604
rect 488540 68552 488592 68604
rect 35164 68484 35216 68536
rect 87144 68484 87196 68536
rect 193956 68484 194008 68536
rect 430580 68484 430632 68536
rect 25504 68416 25556 68468
rect 85764 68416 85816 68468
rect 204444 68416 204496 68468
rect 483020 68416 483072 68468
rect 22744 68348 22796 68400
rect 85120 68348 85172 68400
rect 213552 68348 213604 68400
rect 500960 68348 501012 68400
rect 50988 68280 51040 68332
rect 111800 68280 111852 68332
rect 134524 68280 134576 68332
rect 312544 68280 312596 68332
rect 314752 68280 314804 68332
rect 315304 68280 315356 68332
rect 404268 68280 404320 68332
rect 579620 68280 579672 68332
=======
rect 134524 68552 134576 68604
rect 312544 68552 312596 68604
rect 314752 68552 314804 68604
rect 315304 68552 315356 68604
rect 403716 68552 403768 68604
rect 579620 68552 579672 68604
rect 35164 68484 35216 68536
rect 87144 68484 87196 68536
rect 177304 68484 177356 68536
rect 229560 68484 229612 68536
rect 244372 68484 244424 68536
rect 245568 68484 245620 68536
rect 295984 68484 296036 68536
rect 488540 68484 488592 68536
rect 25504 68416 25556 68468
rect 85764 68416 85816 68468
rect 193956 68416 194008 68468
rect 430580 68416 430632 68468
rect 22744 68348 22796 68400
rect 85120 68348 85172 68400
rect 204444 68348 204496 68400
rect 483020 68348 483072 68400
rect 50988 68280 51040 68332
rect 111800 68280 111852 68332
rect 213644 68280 213696 68332
rect 500960 68280 501012 68332
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 274364 67260 274416 67312
rect 374000 67260 374052 67312
rect 385132 67260 385184 67312
rect 496820 67260 496872 67312
rect 209044 67192 209096 67244
rect 326528 67192 326580 67244
rect 387248 67192 387300 67244
rect 506480 67192 506532 67244
rect 310152 67124 310204 67176
rect 484400 67124 484452 67176
rect 43444 67056 43496 67108
rect 89812 67056 89864 67108
rect 292396 67056 292448 67108
rect 466460 67056 466512 67108
rect 39304 66988 39356 67040
rect 88524 66988 88576 67040
rect 192576 66988 192628 67040
rect 423680 66988 423732 67040
rect 32404 66920 32456 66972
rect 86500 66920 86552 66972
rect 205824 66920 205876 66972
rect 489920 66920 489972 66972
rect 15844 66852 15896 66904
rect 107384 66852 107436 66904
rect 209320 66852 209372 66904
rect 507860 66852 507912 66904
rect 387984 65832 388036 65884
rect 510620 65832 510672 65884
<<<<<<< HEAD
rect 392400 65764 392452 65816
=======
rect 391940 65764 391992 65816
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 524420 65764 524472 65816
rect 289544 65696 289596 65748
rect 463700 65696 463752 65748
rect 82360 65628 82412 65680
rect 114652 65628 114704 65680
rect 293776 65628 293828 65680
rect 470600 65628 470652 65680
rect 197452 65560 197504 65612
rect 448520 65560 448572 65612
rect 53656 65492 53708 65544
rect 115112 65492 115164 65544
rect 222568 65492 222620 65544
rect 575480 65492 575532 65544
rect 383476 64336 383528 64388
rect 485780 64336 485832 64388
rect 390376 64268 390428 64320
rect 517520 64268 517572 64320
rect 394516 64200 394568 64252
rect 539600 64200 539652 64252
rect 288256 64132 288308 64184
rect 456892 64132 456944 64184
rect 393136 62840 393188 62892
rect 530584 62840 530636 62892
rect 395896 62772 395948 62824
rect 546500 62772 546552 62824
rect 406752 60664 406804 60716
rect 580172 60664 580224 60716
rect 389088 58624 389140 58676
rect 514760 58624 514812 58676
rect 235908 50328 235960 50380
rect 331864 50328 331916 50380
rect 394608 50328 394660 50380
rect 542360 50328 542412 50380
rect 45376 48968 45428 49020
rect 87604 48968 87656 49020
rect 176476 48968 176528 49020
rect 338304 48968 338356 49020
rect 175096 47540 175148 47592
rect 331312 47540 331364 47592
rect 406660 46860 406712 46912
rect 580172 46860 580224 46912
rect 228456 44820 228508 44872
rect 328552 44820 328604 44872
rect 406568 33056 406620 33108
rect 579896 33056 579948 33108
rect 238024 25508 238076 25560
rect 331404 25508 331456 25560
rect 289728 24080 289780 24132
rect 459560 24080 459612 24132
rect 227076 22720 227128 22772
rect 329932 22720 329984 22772
rect 393228 22720 393280 22772
rect 535460 22720 535512 22772
rect 268936 21360 268988 21412
rect 354036 21360 354088 21412
rect 390468 21360 390520 21412
rect 521660 21360 521712 21412
rect 406476 20612 406528 20664
rect 579896 20612 579948 20664
rect 295984 19932 296036 19984
rect 342352 19932 342404 19984
rect 198556 18776 198608 18828
rect 236092 18776 236144 18828
rect 222936 18708 222988 18760
rect 329840 18708 329892 18760
rect 202604 18640 202656 18692
rect 327172 18640 327224 18692
rect 162124 18572 162176 18624
rect 313280 18572 313332 18624
rect 386328 18572 386380 18624
rect 499580 18572 499632 18624
rect 249064 17892 249116 17944
rect 251180 17892 251232 17944
rect 242256 17552 242308 17604
rect 334072 17552 334124 17604
rect 271696 17484 271748 17536
rect 367100 17484 367152 17536
rect 177856 17416 177908 17468
rect 231952 17416 232004 17468
rect 232596 17416 232648 17468
rect 328460 17416 328512 17468
rect 195244 17348 195296 17400
rect 324412 17348 324464 17400
rect 178684 17280 178736 17332
rect 320364 17280 320416 17332
rect 175096 17212 175148 17264
rect 321652 17212 321704 17264
rect 383568 17212 383620 17264
rect 481732 17212 481784 17264
rect 270316 16328 270368 16380
rect 354128 16328 354180 16380
rect 271788 16260 271840 16312
<<<<<<< HEAD
rect 371700 16260 371752 16312
=======
rect 371240 16260 371292 16312
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 224408 16192 224460 16244
rect 327080 16192 327132 16244
rect 196624 16124 196676 16176
rect 323124 16124 323176 16176
rect 173256 16056 173308 16108
rect 313464 16056 313516 16108
rect 173164 15988 173216 16040
rect 316316 15988 316368 16040
rect 164148 15920 164200 15972
rect 309784 15920 309836 15972
rect 197176 15852 197228 15904
rect 441528 15852 441580 15904
rect 267556 14968 267608 15020
rect 349344 14968 349396 15020
rect 231216 14900 231268 14952
rect 331220 14900 331272 14952
rect 206376 14832 206428 14884
rect 324320 14832 324372 14884
rect 195336 14764 195388 14816
rect 321560 14764 321612 14816
rect 170956 14696 171008 14748
<<<<<<< HEAD
rect 310244 14696 310296 14748
rect 175188 14628 175240 14680
rect 335084 14628 335136 14680
=======
rect 309784 14696 309836 14748
rect 175188 14628 175240 14680
rect 334624 14628 334676 14680
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 179236 14560 179288 14612
rect 352840 14560 352892 14612
rect 170404 14492 170456 14544
rect 230572 14492 230624 14544
rect 292488 14492 292540 14544
rect 478144 14492 478196 14544
rect 30104 14424 30156 14476
rect 64972 14424 65024 14476
rect 195796 14424 195848 14476
<<<<<<< HEAD
rect 437940 14424 437992 14476
=======
rect 437480 14424 437532 14476
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 104164 14084 104216 14136
rect 105728 14084 105780 14136
rect 173624 13676 173676 13728
rect 231860 13676 231912 13728
rect 270408 13676 270460 13728
rect 360844 13676 360896 13728
rect 195612 13608 195664 13660
rect 287704 13608 287756 13660
rect 231768 13540 231820 13592
rect 327724 13540 327776 13592
rect 169576 13472 169628 13524
<<<<<<< HEAD
rect 306748 13472 306800 13524
=======
rect 306380 13472 306432 13524
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 173808 13404 173860 13456
rect 324412 13404 324464 13456
rect 173716 13336 173768 13388
rect 328000 13336 328052 13388
rect 177764 13268 177816 13320
rect 349252 13268 349304 13320
rect 195888 13200 195940 13252
<<<<<<< HEAD
rect 434444 13200 434496 13252
rect 198648 13132 198700 13184
rect 452108 13132 452160 13184
=======
rect 433984 13200 434036 13252
rect 198648 13132 198700 13184
rect 451648 13132 451700 13184
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 206928 13064 206980 13116
rect 494704 13064 494756 13116
rect 267648 12384 267700 12436
rect 346952 12384 347004 12436
rect 181904 12316 181956 12368
rect 291844 12316 291896 12368
rect 169668 12248 169720 12300
rect 303160 12248 303212 12300
rect 171048 12180 171100 12232
rect 313832 12180 313884 12232
rect 169576 12112 169628 12164
rect 230480 12112 230532 12164
rect 286876 12112 286928 12164
<<<<<<< HEAD
rect 446220 12112 446272 12164
=======
rect 445760 12112 445812 12164
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 160744 12044 160796 12096
rect 227812 12044 227864 12096
rect 286968 12044 287020 12096
rect 449808 12044 449860 12096
rect 162676 11976 162728 12028
rect 267740 11976 267792 12028
rect 288348 11976 288400 12028
rect 453304 11976 453356 12028
rect 176568 11908 176620 11960
rect 341064 11908 341116 11960
rect 353944 11908 353996 11960
<<<<<<< HEAD
rect 427268 11908 427320 11960
rect 165528 11840 165580 11892
rect 285404 11840 285456 11892
rect 296628 11840 296680 11892
rect 499396 11840 499448 11892
=======
rect 426808 11908 426860 11960
rect 165528 11840 165580 11892
rect 284944 11840 284996 11892
rect 296628 11840 296680 11892
rect 498936 11840 498988 11892
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 197268 11772 197320 11824
rect 445024 11772 445076 11824
rect 224316 11704 224368 11756
rect 498200 11704 498252 11756
rect 226984 11636 227036 11688
<<<<<<< HEAD
rect 281908 11636 281960 11688
=======
rect 281540 11636 281592 11688
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 278688 10956 278740 11008
rect 407212 10956 407264 11008
rect 202512 10888 202564 10940
rect 237472 10888 237524 10940
rect 279976 10888 280028 10940
rect 410800 10888 410852 10940
rect 191564 10820 191616 10872
rect 234712 10820 234764 10872
rect 280068 10820 280120 10872
rect 414296 10820 414348 10872
rect 414664 10820 414716 10872
rect 490012 10820 490064 10872
rect 187332 10752 187384 10804
rect 232504 10752 232556 10804
rect 281356 10752 281408 10804
<<<<<<< HEAD
rect 417884 10752 417936 10804
rect 209136 10684 209188 10736
rect 274824 10684 274876 10736
rect 281264 10684 281316 10736
rect 421380 10684 421432 10736
=======
rect 417424 10752 417476 10804
rect 209136 10684 209188 10736
rect 274824 10684 274876 10736
rect 281264 10684 281316 10736
rect 420920 10684 420972 10736
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 162492 10616 162544 10668
rect 228364 10616 228416 10668
rect 282736 10616 282788 10668
rect 424968 10616 425020 10668
rect 158628 10548 158680 10600
rect 249984 10548 250036 10600
rect 250444 10548 250496 10600
rect 278320 10548 278372 10600
rect 282828 10548 282880 10600
rect 428464 10548 428516 10600
rect 159916 10480 159968 10532
rect 253480 10480 253532 10532
rect 284208 10480 284260 10532
rect 432052 10480 432104 10532
rect 161388 10412 161440 10464
<<<<<<< HEAD
rect 259460 10412 259512 10464
rect 284116 10412 284168 10464
rect 435548 10412 435600 10464
=======
rect 260656 10412 260708 10464
rect 284116 10412 284168 10464
rect 435088 10412 435140 10464
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 161296 10344 161348 10396
rect 264152 10344 264204 10396
rect 285496 10344 285548 10396
rect 439136 10344 439188 10396
rect 162768 10276 162820 10328
<<<<<<< HEAD
rect 271236 10276 271288 10328
=======
rect 270776 10276 270828 10328
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 285588 10276 285640 10328
rect 442632 10276 442684 10328
rect 278596 10208 278648 10260
rect 403624 10208 403676 10260
rect 277308 10140 277360 10192
rect 398840 10140 398892 10192
rect 277216 10072 277268 10124
<<<<<<< HEAD
rect 396540 10072 396592 10124
rect 275928 10004 275980 10056
rect 393044 10004 393096 10056
=======
rect 396080 10072 396132 10124
rect 275928 10004 275980 10056
rect 392584 10004 392636 10056
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 275836 9936 275888 9988
rect 389456 9936 389508 9988
rect 274548 9868 274600 9920
rect 385960 9868 386012 9920
rect 274456 9800 274508 9852
rect 382372 9800 382424 9852
rect 273168 9732 273220 9784
<<<<<<< HEAD
rect 378876 9732 378928 9784
=======
rect 378416 9732 378468 9784
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 215668 9596 215720 9648
rect 240232 9596 240284 9648
rect 240508 9596 240560 9648
rect 244372 9596 244424 9648
rect 308956 9596 309008 9648
rect 563244 9596 563296 9648
rect 199936 9528 199988 9580
rect 455696 9528 455748 9580
rect 180248 9460 180300 9512
rect 222844 9460 222896 9512
rect 259276 9460 259328 9512
rect 304356 9460 304408 9512
rect 311808 9460 311860 9512
rect 570328 9460 570380 9512
rect 200028 9392 200080 9444
rect 459192 9392 459244 9444
rect 201408 9324 201460 9376
rect 462780 9324 462832 9376
rect 183744 9256 183796 9308
rect 233332 9256 233384 9308
rect 259368 9256 259420 9308
rect 307944 9256 307996 9308
rect 311716 9256 311768 9308
rect 573916 9256 573968 9308
<<<<<<< HEAD
rect 129648 9188 129700 9240
=======
rect 129556 9188 129608 9240
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 222200 9188 222252 9240
rect 222752 9188 222804 9240
rect 241612 9188 241664 9240
rect 249616 9188 249668 9240
rect 258264 9188 258316 9240
rect 260748 9188 260800 9240
rect 311440 9188 311492 9240
rect 313096 9188 313148 9240
rect 577412 9188 577464 9240
rect 201316 9120 201368 9172
rect 466276 9120 466328 9172
rect 80888 9052 80940 9104
rect 98092 9052 98144 9104
rect 202788 9052 202840 9104
rect 469864 9052 469916 9104
rect 202696 8984 202748 9036
rect 473452 8984 473504 9036
rect 81348 8916 81400 8968
rect 104532 8916 104584 8968
rect 204168 8916 204220 8968
rect 476948 8916 477000 8968
rect 266268 8848 266320 8900
rect 339868 8848 339920 8900
rect 264796 8780 264848 8832
rect 336280 8780 336332 8832
rect 264888 8712 264940 8764
rect 332692 8712 332744 8764
rect 263508 8644 263560 8696
rect 329196 8644 329248 8696
rect 263416 8576 263468 8628
rect 325608 8576 325660 8628
rect 262128 8508 262180 8560
rect 322112 8508 322164 8560
rect 262036 8440 262088 8492
rect 318524 8440 318576 8492
<<<<<<< HEAD
rect 260656 8372 260708 8424
=======
rect 260564 8372 260616 8424
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 315028 8372 315080 8424
rect 184756 8236 184808 8288
rect 384764 8236 384816 8288
rect 186228 8168 186280 8220
rect 388260 8168 388312 8220
rect 187608 8100 187660 8152
rect 391848 8100 391900 8152
rect 187516 8032 187568 8084
rect 395344 8032 395396 8084
rect 188896 7964 188948 8016
rect 398932 7964 398984 8016
rect 188988 7896 189040 7948
rect 402520 7896 402572 7948
rect 190276 7828 190328 7880
rect 406016 7828 406068 7880
rect 411904 7828 411956 7880
rect 480536 7828 480588 7880
rect 190368 7760 190420 7812
rect 409604 7760 409656 7812
rect 410524 7760 410576 7812
rect 495900 7760 495952 7812
rect 191656 7692 191708 7744
rect 413100 7692 413152 7744
rect 413284 7692 413336 7744
rect 505376 7692 505428 7744
rect 83464 7624 83516 7676
rect 93860 7624 93912 7676
rect 191748 7624 191800 7676
rect 416688 7624 416740 7676
rect 418804 7624 418856 7676
rect 492312 7624 492364 7676
rect 51356 7556 51408 7608
rect 69204 7556 69256 7608
rect 70308 7556 70360 7608
rect 94596 7556 94648 7608
rect 106096 7556 106148 7608
rect 116400 7556 116452 7608
rect 193128 7556 193180 7608
rect 420184 7556 420236 7608
rect 184848 7488 184900 7540
rect 381176 7488 381228 7540
rect 183468 7420 183520 7472
rect 377680 7420 377732 7472
rect 183376 7352 183428 7404
rect 374092 7352 374144 7404
rect 181996 7284 182048 7336
rect 370596 7284 370648 7336
rect 371884 7284 371936 7336
rect 487620 7284 487672 7336
rect 182088 7216 182140 7268
rect 367008 7216 367060 7268
rect 180708 7148 180760 7200
rect 363512 7148 363564 7200
rect 180616 7080 180668 7132
rect 359924 7080 359976 7132
rect 179328 7012 179380 7064
rect 356336 7012 356388 7064
rect 206284 6808 206336 6860
rect 232228 6808 232280 6860
rect 255228 6808 255280 6860
rect 283104 6808 283156 6860
rect 302056 6808 302108 6860
rect 527824 6808 527876 6860
rect 205088 6740 205140 6792
rect 237380 6740 237432 6792
rect 255136 6740 255188 6792
rect 286600 6740 286652 6792
rect 303528 6740 303580 6792
rect 531320 6740 531372 6792
rect 204904 6672 204956 6724
rect 239312 6672 239364 6724
rect 256608 6672 256660 6724
rect 290188 6672 290240 6724
rect 303436 6672 303488 6724
rect 534908 6672 534960 6724
rect 155776 6604 155828 6656
rect 235816 6604 235868 6656
rect 237012 6604 237064 6656
rect 244280 6604 244332 6656
rect 256516 6604 256568 6656
rect 293684 6604 293736 6656
rect 304816 6604 304868 6656
rect 538404 6604 538456 6656
rect 157248 6536 157300 6588
rect 242900 6536 242952 6588
rect 257896 6536 257948 6588
rect 297272 6536 297324 6588
rect 304908 6536 304960 6588
rect 541992 6536 542044 6588
rect 79324 6468 79376 6520
rect 90364 6468 90416 6520
rect 160008 6468 160060 6520
rect 257068 6468 257120 6520
rect 257988 6468 258040 6520
rect 300768 6468 300820 6520
rect 306196 6468 306248 6520
rect 545488 6468 545540 6520
rect 167184 6400 167236 6452
rect 289084 6400 289136 6452
rect 306288 6400 306340 6452
rect 549076 6400 549128 6452
rect 42800 6332 42852 6384
rect 89904 6332 89956 6384
rect 166816 6332 166868 6384
rect 288992 6332 289044 6384
rect 307668 6332 307720 6384
rect 552664 6332 552716 6384
rect 34796 6264 34848 6316
rect 88340 6264 88392 6316
rect 166908 6264 166960 6316
rect 292580 6264 292632 6316
rect 307576 6264 307628 6316
rect 556160 6264 556212 6316
rect 2872 6196 2924 6248
rect 57244 6196 57296 6248
rect 63224 6196 63276 6248
rect 93952 6196 94004 6248
rect 168288 6196 168340 6248
rect 296076 6196 296128 6248
rect 309048 6196 309100 6248
rect 559748 6196 559800 6248
rect 27712 6128 27764 6180
rect 86960 6128 87012 6180
rect 87972 6128 88024 6180
rect 98644 6128 98696 6180
rect 141884 6128 141936 6180
rect 164884 6128 164936 6180
rect 168196 6128 168248 6180
rect 299664 6128 299716 6180
rect 310428 6128 310480 6180
rect 566832 6128 566884 6180
rect 204996 6060 205048 6112
rect 228732 6060 228784 6112
rect 229836 6060 229888 6112
rect 242164 6060 242216 6112
rect 253756 6060 253808 6112
rect 279516 6060 279568 6112
rect 302148 6060 302200 6112
rect 524236 6060 524288 6112
rect 224224 5992 224276 6044
rect 246396 5992 246448 6044
rect 253848 5992 253900 6044
rect 276020 5992 276072 6044
rect 300676 5992 300728 6044
rect 520740 5992 520792 6044
rect 219256 5924 219308 5976
rect 240140 5924 240192 5976
rect 252376 5924 252428 5976
rect 272432 5924 272484 5976
rect 300584 5924 300636 5976
rect 517152 5924 517204 5976
rect 212172 5856 212224 5908
rect 231124 5856 231176 5908
rect 251088 5856 251140 5908
rect 261760 5856 261812 5908
rect 299204 5856 299256 5908
rect 513564 5856 513616 5908
rect 299296 5788 299348 5840
rect 510068 5788 510120 5840
rect 297916 5720 297968 5772
<<<<<<< HEAD
rect 506572 5720 506624 5772
=======
rect 506480 5720 506532 5772
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 298008 5652 298060 5704
rect 502984 5652 503036 5704
rect 406384 5584 406436 5636
rect 580172 5584 580224 5636
rect 69112 5516 69164 5568
rect 72424 5516 72476 5568
rect 98644 5516 98696 5568
rect 100760 5516 100812 5568
rect 104716 5516 104768 5568
rect 112812 5516 112864 5568
rect 244096 5516 244148 5568
rect 245660 5516 245712 5568
rect 246948 5516 247000 5568
rect 247592 5516 247644 5568
rect 249708 5516 249760 5568
rect 254676 5516 254728 5568
rect 146208 5448 146260 5500
rect 186136 5448 186188 5500
rect 215208 5448 215260 5500
rect 537208 5448 537260 5500
rect 79968 5380 80020 5432
rect 97448 5380 97500 5432
rect 147588 5380 147640 5432
rect 189724 5380 189776 5432
rect 216496 5380 216548 5432
rect 540796 5380 540848 5432
rect 84476 5312 84528 5364
rect 98000 5312 98052 5364
rect 147496 5312 147548 5364
rect 193220 5312 193272 5364
rect 216588 5312 216640 5364
rect 544384 5312 544436 5364
rect 77392 5244 77444 5296
rect 96804 5244 96856 5296
rect 148876 5244 148928 5296
rect 196808 5244 196860 5296
rect 217876 5244 217928 5296
rect 547880 5244 547932 5296
rect 79876 5176 79928 5228
rect 101036 5176 101088 5228
rect 148784 5176 148836 5228
rect 200304 5176 200356 5228
rect 217968 5176 218020 5228
rect 551468 5176 551520 5228
rect 52552 5108 52604 5160
rect 65524 5108 65576 5160
rect 73804 5108 73856 5160
rect 96712 5108 96764 5160
rect 150256 5108 150308 5160
rect 203892 5108 203944 5160
rect 219164 5108 219216 5160
rect 554964 5108 555016 5160
rect 44272 5040 44324 5092
rect 67732 5040 67784 5092
rect 77208 5040 77260 5092
rect 85764 5040 85816 5092
rect 86224 5040 86276 5092
rect 111616 5040 111668 5092
rect 150348 5040 150400 5092
rect 207388 5040 207440 5092
rect 219348 5040 219400 5092
rect 558552 5040 558604 5092
rect 21824 4972 21876 5024
rect 53104 4972 53156 5024
rect 59636 4972 59688 5024
rect 93124 4972 93176 5024
rect 151728 4972 151780 5024
rect 210976 4972 211028 5024
rect 220636 4972 220688 5024
rect 562048 4972 562100 5024
rect 4068 4904 4120 4956
rect 50344 4904 50396 4956
rect 56048 4904 56100 4956
rect 92572 4904 92624 4956
rect 106188 4904 106240 4956
rect 116492 4904 116544 4956
rect 151636 4904 151688 4956
rect 214472 4904 214524 4956
rect 220728 4904 220780 4956
rect 565636 4904 565688 4956
rect 7656 4836 7708 4888
rect 60832 4836 60884 4888
rect 62028 4836 62080 4888
rect 69664 4836 69716 4888
rect 84108 4836 84160 4888
rect 118792 4836 118844 4888
rect 153016 4836 153068 4888
rect 218060 4836 218112 4888
rect 222108 4836 222160 4888
rect 569132 4836 569184 4888
rect 572 4768 624 4820
rect 58624 4768 58676 4820
rect 84016 4768 84068 4820
rect 122288 4768 122340 4820
rect 153108 4768 153160 4820
rect 221556 4768 221608 4820
rect 222016 4768 222068 4820
rect 572720 4768 572772 4820
rect 58440 4700 58492 4752
rect 70584 4700 70636 4752
rect 146116 4700 146168 4752
rect 182548 4700 182600 4752
rect 215116 4700 215168 4752
rect 533712 4700 533764 4752
rect 144644 4632 144696 4684
rect 179052 4632 179104 4684
rect 213736 4632 213788 4684
rect 530124 4632 530176 4684
rect 144552 4564 144604 4616
rect 175464 4564 175516 4616
rect 213828 4564 213880 4616
rect 526628 4564 526680 4616
rect 91560 4496 91612 4548
rect 94504 4496 94556 4548
rect 143356 4496 143408 4548
rect 171968 4496 172020 4548
rect 212448 4496 212500 4548
rect 523040 4496 523092 4548
rect 143448 4428 143500 4480
rect 168380 4428 168432 4480
rect 212356 4428 212408 4480
rect 519544 4428 519596 4480
rect 211068 4360 211120 4412
rect 515956 4360 516008 4412
rect 210884 4292 210936 4344
rect 512460 4292 512512 4344
rect 65524 4224 65576 4276
rect 71964 4224 72016 4276
rect 75828 4224 75880 4276
rect 79692 4224 79744 4276
<<<<<<< HEAD
rect 109224 4224 109276 4276
rect 154488 4224 154540 4276
rect 225144 4224 225196 4276
=======
rect 154488 4224 154540 4276
rect 225144 4224 225196 4276
rect 252468 4224 252520 4276
rect 268844 4224 268896 4276
rect 269028 4224 269080 4276
rect 354036 4224 354088 4276
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 48964 4156 49016 4208
rect 51724 4156 51776 4208
rect 66720 4156 66772 4208
rect 68284 4156 68336 4208
rect 75736 4156 75788 4208
rect 76196 4156 76248 4208
rect 77116 4156 77168 4208
rect 83280 4156 83332 4208
rect 85764 4156 85816 4208
rect 86868 4156 86920 4208
rect 95148 4156 95200 4208
rect 100944 4156 100996 4208
rect 104808 4156 104860 4208
rect 109316 4156 109368 4208
rect 194416 4156 194468 4208
rect 198004 4156 198056 4208
<<<<<<< HEAD
rect 252468 4156 252520 4208
rect 268844 4224 268896 4276
rect 269028 4224 269080 4276
rect 354036 4224 354088 4276
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 472624 4156 472676 4208
rect 474556 4156 474608 4208
rect 64328 4088 64380 4140
rect 116032 4088 116084 4140
<<<<<<< HEAD
rect 137744 4088 137796 4140
rect 143540 4088 143592 4140
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 266544 4088 266596 4140
rect 339592 4088 339644 4140
rect 361396 4088 361448 4140
rect 372896 4088 372948 4140
rect 379428 4088 379480 4140
rect 465172 4088 465224 4140
rect 60832 4020 60884 4072
rect 116124 4020 116176 4072
rect 216864 4020 216916 4072
rect 227076 4020 227128 4072
rect 262956 4020 263008 4072
rect 338120 4020 338172 4072
<<<<<<< HEAD
rect 344560 4020 344612 4072
rect 354680 4020 354732 4072
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 380808 4020 380860 4072
rect 472256 4020 472308 4072
rect 14740 3952 14792 4004
rect 18604 3952 18656 4004
rect 57244 3952 57296 4004
<<<<<<< HEAD
rect 107752 3952 107804 4004
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 188528 3952 188580 4004
rect 195244 3952 195296 4004
rect 223948 3952 224000 4004
rect 238024 3952 238076 4004
<<<<<<< HEAD
rect 259552 3952 259604 4004
rect 338396 3952 338448 4004
=======
rect 259460 3952 259512 4004
rect 338396 3952 338448 4004
rect 344560 3952 344612 4004
rect 354680 3952 354732 4004
rect 361488 3952 361540 4004
rect 376484 3952 376536 4004
rect 382188 3952 382240 4004
rect 479340 3952 479392 4004
rect 489920 3952 489972 4004
rect 491116 3952 491168 4004
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 46664 3884 46716 3936
rect 31300 3816 31352 3868
rect 39304 3816 39356 3868
rect 43076 3816 43128 3868
rect 111984 3816 112036 3868
rect 23020 3748 23072 3800
rect 35164 3748 35216 3800
rect 39580 3748 39632 3800
rect 111892 3748 111944 3800
rect 25504 3680 25556 3732
rect 38384 3680 38436 3732
rect 43444 3680 43496 3732
rect 110604 3680 110656 3732
rect 15936 3612 15988 3664
rect 21364 3612 21416 3664
rect 6460 3544 6512 3596
rect 11704 3544 11756 3596
rect 13544 3544 13596 3596
rect 9956 3476 10008 3528
rect 15844 3476 15896 3528
rect 22744 3544 22796 3596
rect 1676 3408 1728 3460
rect 7564 3408 7616 3460
rect 8760 3408 8812 3460
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 18236 3476 18288 3528
rect 32312 3612 32364 3664
rect 32404 3612 32456 3664
rect 110512 3612 110564 3664
rect 28908 3544 28960 3596
rect 109132 3544 109184 3596
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 24216 3408 24268 3460
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
<<<<<<< HEAD
=======
rect 109224 3476 109276 3528
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 110512 3476 110564 3528
rect 111708 3476 111760 3528
rect 140596 3884 140648 3936
rect 157800 3884 157852 3936
rect 158904 3884 158956 3936
rect 177304 3884 177356 3936
rect 192024 3884 192076 3936
rect 206376 3884 206428 3936
rect 209780 3884 209832 3936
rect 131764 3816 131816 3868
rect 162124 3816 162176 3868
rect 170772 3816 170824 3868
rect 178684 3816 178736 3868
rect 184940 3816 184992 3868
rect 196624 3816 196676 3868
rect 206192 3816 206244 3868
rect 224408 3816 224460 3868
rect 227536 3884 227588 3936
rect 231216 3884 231268 3936
rect 255872 3884 255924 3936
rect 336832 3884 336884 3936
rect 228456 3816 228508 3868
rect 252376 3816 252428 3868
rect 336740 3816 336792 3868
<<<<<<< HEAD
rect 341156 3816 341208 3868
=======
rect 340972 3816 341024 3868
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 135260 3748 135312 3800
rect 173256 3748 173308 3800
rect 177948 3748 178000 3800
rect 195336 3748 195388 3800
rect 199108 3748 199160 3800
rect 209044 3748 209096 3800
rect 213368 3748 213420 3800
rect 232596 3748 232648 3800
rect 238116 3748 238168 3800
rect 242256 3748 242308 3800
rect 248788 3748 248840 3800
rect 335452 3748 335504 3800
<<<<<<< HEAD
rect 340972 3748 341024 3800
rect 342076 3748 342128 3800
rect 142068 3680 142120 3732
rect 160100 3680 160152 3732
rect 316132 3680 316184 3732
rect 316408 3680 316460 3732
rect 333888 3680 333940 3732
rect 352012 3952 352064 4004
rect 361488 3952 361540 4004
rect 376484 3952 376536 4004
rect 382188 3952 382240 4004
rect 479340 3952 479392 4004
rect 349436 3927 349488 3936
rect 349436 3893 349445 3927
rect 349445 3893 349479 3927
rect 349479 3893 349488 3927
rect 349436 3884 349488 3893
=======
rect 343732 3748 343784 3800
rect 142068 3680 142120 3732
rect 160100 3680 160152 3732
rect 318892 3680 318944 3732
rect 333888 3680 333940 3732
rect 352012 3884 352064 3936
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 360844 3884 360896 3936
rect 364616 3884 364668 3936
rect 397368 3884 397420 3936
rect 550272 3884 550324 3936
rect 362868 3816 362920 3868
rect 379980 3816 380032 3868
rect 397276 3816 397328 3868
rect 553768 3816 553820 3868
<<<<<<< HEAD
rect 139216 3612 139268 3664
rect 137836 3544 137888 3596
rect 140044 3544 140096 3596
rect 140688 3612 140740 3664
rect 154212 3612 154264 3664
rect 156604 3612 156656 3664
=======
rect 140688 3612 140740 3664
rect 154212 3612 154264 3664
rect 156604 3612 156656 3664
rect 139216 3544 139268 3596
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 150624 3544 150676 3596
rect 153016 3544 153068 3596
rect 317512 3612 317564 3664
rect 319720 3612 319772 3664
rect 312636 3544 312688 3596
rect 313188 3544 313240 3596
rect 316224 3544 316276 3596
rect 113272 3476 113324 3528
<<<<<<< HEAD
rect 118976 3476 119028 3528
=======
rect 114008 3476 114060 3528
rect 114468 3476 114520 3528
rect 121644 3476 121696 3528
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 125876 3476 125928 3528
rect 126888 3476 126940 3528
<<<<<<< HEAD
=======
rect 126980 3476 127032 3528
rect 129556 3476 129608 3528
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 130568 3476 130620 3528
rect 131028 3476 131080 3528
rect 132960 3476 133012 3528
rect 133788 3476 133840 3528
<<<<<<< HEAD
rect 19432 3340 19484 3392
rect 114560 3408 114612 3460
rect 121644 3408 121696 3460
rect 128176 3408 128228 3460
rect 134524 3476 134576 3528
rect 139308 3476 139360 3528
rect 147128 3476 147180 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 149520 3476 149572 3528
rect 317604 3476 317656 3528
rect 134156 3408 134208 3460
rect 135168 3408 135220 3460
rect 145932 3408 145984 3460
rect 316040 3408 316092 3460
rect 316132 3408 316184 3460
rect 318892 3408 318944 3460
rect 323308 3408 323360 3460
rect 324228 3408 324280 3460
=======
rect 141240 3476 141292 3528
rect 141976 3476 142028 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 149520 3476 149572 3528
rect 316408 3476 316460 3528
rect 19432 3340 19484 3392
rect 107844 3408 107896 3460
rect 114560 3408 114612 3460
rect 121552 3408 121604 3460
rect 128176 3408 128228 3460
rect 134524 3408 134576 3460
rect 139308 3408 139360 3460
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 50160 3340 50212 3392
rect 50988 3340 51040 3392
rect 67916 3340 67968 3392
rect 117412 3340 117464 3392
rect 137836 3340 137888 3392
rect 140044 3340 140096 3392
rect 145932 3408 145984 3460
rect 316040 3408 316092 3460
rect 317604 3408 317656 3460
rect 323308 3476 323360 3528
rect 324228 3476 324280 3528
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 330392 3612 330444 3664
rect 351920 3748 351972 3800
rect 362776 3748 362828 3800
rect 383568 3748 383620 3800
rect 395988 3748 396040 3800
rect 399944 3748 399996 3800
rect 557356 3748 557408 3800
rect 364248 3680 364300 3732
rect 387156 3680 387208 3732
rect 398748 3680 398800 3732
rect 560852 3680 560904 3732
rect 326804 3544 326856 3596
rect 350724 3612 350776 3664
rect 353944 3612 353996 3664
rect 357532 3612 357584 3664
rect 360016 3612 360068 3664
rect 348056 3544 348108 3596
rect 354772 3544 354824 3596
rect 358636 3544 358688 3596
rect 362316 3544 362368 3596
rect 364156 3612 364208 3664
rect 390652 3612 390704 3664
rect 398656 3612 398708 3664
rect 564440 3612 564492 3664
rect 369400 3544 369452 3596
rect 349160 3476 349212 3528
rect 355232 3476 355284 3528
rect 356244 3476 356296 3528
rect 357440 3476 357492 3528
rect 358728 3476 358780 3528
rect 365628 3476 365680 3528
rect 394240 3544 394292 3596
rect 400036 3544 400088 3596
rect 568028 3544 568080 3596
<<<<<<< HEAD
=======
rect 349436 3408 349488 3460
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 354128 3408 354180 3460
rect 361120 3408 361172 3460
rect 365536 3408 365588 3460
rect 397736 3476 397788 3528
rect 398840 3476 398892 3528
rect 400128 3476 400180 3528
rect 571524 3476 571576 3528
<<<<<<< HEAD
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 50160 3340 50212 3392
rect 50988 3340 51040 3392
rect 72608 3340 72660 3392
rect 73068 3340 73120 3392
rect 35992 3272 36044 3324
rect 67916 3204 67968 3256
rect 117412 3340 117464 3392
=======
rect 147128 3340 147180 3392
rect 155408 3340 155460 3392
rect 155868 3340 155920 3392
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 161296 3340 161348 3392
rect 163688 3340 163740 3392
rect 164148 3340 164200 3392
rect 173164 3340 173216 3392
rect 173624 3340 173676 3392
rect 174268 3340 174320 3392
rect 175096 3340 175148 3392
rect 176660 3340 176712 3392
rect 177856 3340 177908 3392
rect 181444 3340 181496 3392
rect 181904 3340 181956 3392
<<<<<<< HEAD
rect 197912 3340 197964 3392
rect 198556 3340 198608 3392
=======
rect 190828 3340 190880 3392
rect 191564 3340 191616 3392
rect 197912 3340 197964 3392
rect 198556 3340 198608 3392
rect 201500 3340 201552 3392
rect 202512 3340 202564 3392
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 208584 3340 208636 3392
rect 209688 3340 209740 3392
rect 226340 3340 226392 3392
rect 227628 3340 227680 3392
rect 231032 3340 231084 3392
rect 231768 3340 231820 3392
rect 233424 3340 233476 3392
rect 234528 3340 234580 3392
<<<<<<< HEAD
rect 259460 3340 259512 3392
rect 260656 3340 260708 3392
rect 270040 3340 270092 3392
rect 71504 3136 71556 3188
rect 75000 3204 75052 3256
rect 114008 3272 114060 3324
rect 114468 3272 114520 3324
rect 121552 3272 121604 3324
rect 151820 3272 151872 3324
rect 160744 3272 160796 3324
rect 273628 3272 273680 3324
rect 337476 3340 337528 3392
rect 338028 3340 338080 3392
rect 339684 3272 339736 3324
=======
rect 234620 3340 234672 3392
rect 235908 3340 235960 3392
rect 270040 3340 270092 3392
rect 339684 3340 339736 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 346492 3340 346544 3392
rect 35992 3272 36044 3324
rect 71504 3272 71556 3324
rect 117320 3272 117372 3324
rect 273628 3272 273680 3324
rect 72608 3204 72660 3256
rect 73068 3204 73120 3256
rect 75000 3204 75052 3256
rect 118976 3204 119028 3256
rect 277124 3204 277176 3256
rect 41880 3136 41932 3188
rect 42800 3136 42852 3188
rect 78588 3136 78640 3188
rect 118700 3136 118752 3188
rect 134156 3136 134208 3188
rect 135168 3136 135220 3188
rect 166080 3136 166132 3188
rect 170404 3136 170456 3188
rect 284300 3136 284352 3188
rect 337476 3272 337528 3324
rect 338028 3272 338080 3324
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 366824 3272 366876 3324
rect 401324 3408 401376 3460
rect 401508 3408 401560 3460
rect 575112 3408 575164 3460
rect 378048 3340 378100 3392
rect 458088 3340 458140 3392
<<<<<<< HEAD
rect 489920 3340 489972 3392
rect 491116 3340 491168 3392
rect 506480 3340 506532 3392
rect 507676 3340 507728 3392
rect 530584 3340 530636 3392
rect 532516 3340 532568 3392
rect 375196 3272 375248 3324
rect 117320 3204 117372 3256
rect 277124 3204 277176 3256
rect 340880 3204 340932 3256
=======
rect 530584 3340 530636 3392
rect 532516 3340 532568 3392
rect 375196 3272 375248 3324
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 374000 3204 374052 3256
rect 375288 3204 375340 3256
rect 376668 3272 376720 3324
rect 450912 3272 450964 3324
rect 443828 3204 443880 3256
<<<<<<< HEAD
rect 78588 3136 78640 3188
rect 118700 3136 118752 3188
rect 155408 3136 155460 3188
rect 155868 3136 155920 3188
rect 166080 3136 166132 3188
rect 170404 3136 170456 3188
rect 234620 3136 234672 3188
rect 235908 3136 235960 3188
rect 284300 3136 284352 3188
rect 342444 3136 342496 3188
rect 360108 3136 360160 3188
rect 365812 3136 365864 3188
rect 373908 3136 373960 3188
rect 436744 3136 436796 3188
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 12348 3068 12400 3120
rect 14464 3068 14516 3120
rect 82084 3068 82136 3120
rect 120264 3068 120316 3120
<<<<<<< HEAD
rect 126980 3068 127032 3120
rect 129648 3068 129700 3120
rect 201500 3068 201552 3120
rect 202512 3068 202564 3120
rect 280712 3068 280764 3120
rect 281448 3068 281500 3120
rect 287796 3068 287848 3120
rect 343640 3068 343692 3120
rect 371148 3068 371200 3120
rect 426164 3068 426216 3120
rect 431960 3068 432012 3120
rect 433248 3068 433300 3120
=======
rect 280712 3068 280764 3120
rect 281448 3068 281500 3120
rect 287796 3068 287848 3120
rect 341156 3136 341208 3188
rect 360108 3136 360160 3188
rect 365812 3136 365864 3188
rect 373908 3136 373960 3188
rect 436744 3136 436796 3188
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 85672 3000 85724 3052
rect 89168 2932 89220 2984
rect 117596 3000 117648 3052
rect 119344 3000 119396 3052
<<<<<<< HEAD
rect 141240 3000 141292 3052
rect 141976 3000 142028 3052
rect 120172 2932 120224 2984
rect 291384 2932 291436 2984
rect 343732 3000 343784 3052
=======
rect 137744 3000 137796 3052
rect 143540 3000 143592 3052
rect 120172 2932 120224 2984
rect 151820 2932 151872 2984
rect 160744 2932 160796 2984
rect 291384 2932 291436 2984
rect 342444 3068 342496 3120
rect 371148 3068 371200 3120
rect 426164 3068 426216 3120
rect 431960 3068 432012 3120
rect 433248 3068 433300 3120
rect 343640 3000 343692 3052
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 369768 3000 369820 3052
rect 418988 3000 419040 3052
rect 298468 2932 298520 2984
rect 299388 2932 299440 2984
rect 301964 2932 302016 2984
<<<<<<< HEAD
rect 346400 2932 346452 2984
rect 351644 2932 351696 2984
rect 356152 2932 356204 2984
rect 369676 2932 369728 2984
rect 415492 2932 415544 2984
rect 41880 2864 41932 2916
rect 42800 2864 42852 2916
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 92756 2864 92808 2916
rect 116492 2864 116544 2916
rect 119896 2864 119948 2916
rect 135444 2864 135496 2916
rect 136456 2864 136508 2916
<<<<<<< HEAD
rect 190828 2864 190880 2916
rect 191564 2864 191616 2916
rect 220452 2864 220504 2916
rect 222936 2864 222988 2916
rect 305552 2864 305604 2916
rect 346492 2864 346544 2916
rect 368388 2864 368440 2916
rect 96252 2796 96304 2848
rect 99840 2796 99892 2848
rect 100300 2796 100352 2848
=======
rect 220452 2864 220504 2916
rect 222936 2864 222988 2916
rect 305552 2864 305604 2916
rect 351644 2932 351696 2984
rect 356152 2932 356204 2984
rect 369676 2932 369728 2984
rect 415492 2932 415544 2984
rect 346400 2864 346452 2916
rect 368388 2864 368440 2916
rect 96252 2796 96304 2848
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 122932 2796 122984 2848
rect 309048 2796 309100 2848
rect 347964 2796 348016 2848
rect 366916 2796 366968 2848
rect 404820 2796 404872 2848
rect 407120 2864 407172 2916
rect 408408 2864 408460 2916
rect 411904 2796 411956 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 697368 3478 697377
rect 3422 697303 3478 697312
rect 3146 684312 3202 684321
rect 3146 684247 3202 684256
rect 3160 683194 3188 684247
rect 3148 683188 3200 683194
rect 3148 683130 3200 683136
rect 3146 658200 3202 658209
rect 3146 658135 3202 658144
rect 3160 656946 3188 658135
rect 3148 656940 3200 656946
rect 3148 656882 3200 656888
rect 3332 632120 3384 632126
rect 3330 632088 3332 632097
rect 3384 632088 3386 632097
rect 3330 632023 3386 632032
rect 2962 619168 3018 619177
rect 2962 619103 3018 619112
rect 2976 618322 3004 619103
rect 2964 618316 3016 618322
rect 2964 618258 3016 618264
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 2778 593056 2834 593065
rect 2778 592991 2834 593000
rect 2792 592346 2820 592991
rect 2780 592340 2832 592346
rect 2780 592282 2832 592288
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3330 540832 3386 540841
rect 3330 540767 3386 540776
rect 3344 539714 3372 540767
rect 3332 539708 3384 539714
rect 3332 539650 3384 539656
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3344 527202 3372 527847
rect 3332 527196 3384 527202
rect 3332 527138 3384 527144
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 2870 475688 2926 475697
rect 2870 475623 2926 475632
rect 2884 474774 2912 475623
rect 2872 474768 2924 474774
rect 2872 474710 2924 474716
rect 3054 462632 3110 462641
rect 3054 462567 3110 462576
rect 3068 462398 3096 462567
rect 3056 462392 3108 462398
rect 3056 462334 3108 462340
rect 2962 449576 3018 449585
rect 2962 449511 3018 449520
rect 2976 448594 3004 449511
rect 2964 448588 3016 448594
rect 2964 448530 3016 448536
rect 2962 423600 3018 423609
rect 2962 423535 3018 423544
rect 2976 422346 3004 423535
rect 2964 422340 3016 422346
rect 2964 422282 3016 422288
rect 3330 384432 3386 384441
rect 3330 384367 3386 384376
rect 3238 371376 3294 371385
rect 3238 371311 3294 371320
rect 3146 319288 3202 319297
rect 3146 319223 3202 319232
rect 3054 306232 3110 306241
rect 3054 306167 3110 306176
rect 2962 293176 3018 293185
rect 2962 293111 3018 293120
rect 2870 254144 2926 254153
rect 2870 254079 2926 254088
rect 2884 178022 2912 254079
rect 2976 194546 3004 293111
rect 3068 200122 3096 306167
rect 3160 205630 3188 319223
rect 3252 227730 3280 371311
rect 3344 233238 3372 384367
rect 3436 365702 3464 697303
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3424 365696 3476 365702
rect 3424 365638 3476 365644
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3332 233232 3384 233238
rect 3332 233174 3384 233180
rect 3240 227724 3292 227730
rect 3240 227666 3292 227672
rect 3436 222154 3464 358391
rect 3528 356046 3556 671191
rect 3606 645144 3662 645153
rect 3606 645079 3662 645088
rect 3516 356040 3568 356046
rect 3516 355982 3568 355988
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3424 222148 3476 222154
rect 3424 222090 3476 222096
rect 3528 216646 3556 345335
rect 3620 345030 3648 645079
rect 4804 592340 4856 592346
rect 4804 592282 4856 592288
rect 3698 514856 3754 514865
rect 3698 514791 3754 514800
rect 3608 345024 3660 345030
rect 3608 344966 3660 344972
rect 3606 332344 3662 332353
rect 3606 332279 3662 332288
rect 3516 216640 3568 216646
rect 3516 216582 3568 216588
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3148 205624 3200 205630
rect 3148 205566 3200 205572
rect 3056 200116 3108 200122
rect 3056 200058 3108 200064
rect 2964 194540 3016 194546
rect 2964 194482 3016 194488
rect 2872 178016 2924 178022
rect 2872 177958 2924 177964
rect 3436 161430 3464 214911
rect 3620 211138 3648 332279
rect 3712 288386 3740 514791
rect 3790 488744 3846 488753
rect 3790 488679 3846 488688
rect 3700 288380 3752 288386
rect 3700 288322 3752 288328
rect 3698 280120 3754 280129
rect 3698 280055 3754 280064
rect 3608 211132 3660 211138
rect 3608 211074 3660 211080
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3424 161424 3476 161430
rect 3424 161366 3476 161372
rect 3528 155922 3556 201855
rect 3712 189038 3740 280055
rect 3804 277370 3832 488679
rect 3882 436656 3938 436665
rect 3882 436591 3938 436600
rect 3792 277364 3844 277370
rect 3792 277306 3844 277312
rect 3790 267200 3846 267209
rect 3790 267135 3846 267144
rect 3700 189032 3752 189038
rect 3700 188974 3752 188980
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 3516 155916 3568 155922
rect 3516 155858 3568 155864
rect 3620 150414 3648 188799
rect 3804 183530 3832 267135
rect 3896 255270 3924 436591
rect 3974 410544 4030 410553
rect 3974 410479 4030 410488
rect 3884 255264 3936 255270
rect 3884 255206 3936 255212
rect 3988 244254 4016 410479
rect 4066 397488 4122 397497
rect 4066 397423 4122 397432
rect 3976 244248 4028 244254
rect 3976 244190 4028 244196
rect 3882 241088 3938 241097
rect 3882 241023 3938 241032
rect 3792 183524 3844 183530
rect 3792 183466 3844 183472
rect 3698 175944 3754 175953
rect 3698 175879 3754 175888
rect 3608 150408 3660 150414
rect 3608 150350 3660 150356
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3436 133890 3464 149767
rect 3712 144906 3740 175879
rect 3896 172514 3924 241023
rect 4080 238746 4108 397423
rect 4816 322930 4844 592282
rect 7564 539708 7616 539714
rect 7564 539650 7616 539656
rect 4804 322924 4856 322930
rect 4804 322866 4856 322872
rect 7576 299470 7604 539650
rect 8220 369170 8248 702406
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 56796 700398 56824 703520
rect 72988 702434 73016 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 72988 702406 73108 702434
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 56784 700392 56836 700398
rect 56784 700334 56836 700340
rect 71044 700392 71096 700398
rect 71044 700334 71096 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 11704 683188 11756 683194
rect 11704 683130 11756 683136
rect 8208 369164 8260 369170
rect 8208 369106 8260 369112
rect 11716 361554 11744 683130
rect 22744 656940 22796 656946
rect 22744 656882 22796 656888
rect 14464 632120 14516 632126
rect 14464 632062 14516 632068
rect 11704 361548 11756 361554
rect 11704 361490 11756 361496
rect 14476 339454 14504 632062
rect 15844 579692 15896 579698
rect 15844 579634 15896 579640
rect 14464 339448 14516 339454
rect 14464 339390 14516 339396
rect 15856 317422 15884 579634
rect 17224 527196 17276 527202
rect 17224 527138 17276 527144
rect 15844 317416 15896 317422
rect 15844 317358 15896 317364
rect 7564 299464 7616 299470
rect 7564 299406 7616 299412
rect 17236 293962 17264 527138
rect 18604 474768 18656 474774
rect 18604 474710 18656 474716
rect 17224 293956 17276 293962
rect 17224 293898 17276 293904
rect 18616 271862 18644 474710
rect 21364 422340 21416 422346
rect 21364 422282 21416 422288
rect 18604 271856 18656 271862
rect 18604 271798 18656 271804
rect 21376 249762 21404 422282
rect 22756 350538 22784 656882
rect 24780 369238 24808 699654
rect 35164 618316 35216 618322
rect 35164 618258 35216 618264
rect 25504 605872 25556 605878
rect 25504 605814 25556 605820
rect 24768 369232 24820 369238
rect 24768 369174 24820 369180
rect 22744 350532 22796 350538
rect 22744 350474 22796 350480
rect 25516 328438 25544 605814
rect 29644 553444 29696 553450
rect 29644 553386 29696 553392
rect 25504 328432 25556 328438
rect 25504 328374 25556 328380
rect 29656 304978 29684 553386
rect 32404 501016 32456 501022
rect 32404 500958 32456 500964
rect 29644 304972 29696 304978
rect 29644 304914 29696 304920
rect 32416 282878 32444 500958
rect 33784 448588 33836 448594
rect 33784 448530 33836 448536
rect 32404 282872 32456 282878
rect 32404 282814 32456 282820
rect 33796 260846 33824 448530
rect 35176 333946 35204 618258
rect 36544 565888 36596 565894
rect 36544 565830 36596 565836
rect 35164 333940 35216 333946
rect 35164 333882 35216 333888
rect 36556 310486 36584 565830
rect 39304 462392 39356 462398
rect 39304 462334 39356 462340
rect 36544 310480 36596 310486
rect 36544 310422 36596 310428
rect 39316 266354 39344 462334
rect 41340 369306 41368 700334
rect 62028 700324 62080 700330
rect 62028 700266 62080 700272
rect 62040 369850 62068 700266
rect 60832 369844 60884 369850
rect 60832 369786 60884 369792
rect 62028 369844 62080 369850
rect 62028 369786 62080 369792
rect 41328 369300 41380 369306
rect 41328 369242 41380 369248
rect 60844 366194 60872 369786
rect 71056 369374 71084 700334
rect 71044 369368 71096 369374
rect 71044 369310 71096 369316
rect 73080 369170 73108 702406
rect 89444 369300 89496 369306
rect 89444 369242 89496 369248
rect 79600 369232 79652 369238
rect 79600 369174 79652 369180
rect 69756 369164 69808 369170
rect 69756 369106 69808 369112
rect 73068 369164 73120 369170
rect 73068 369106 73120 369112
rect 69768 366194 69796 369106
rect 79612 366194 79640 369174
rect 89456 366194 89484 369242
rect 89640 369238 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 105464 699718 105492 703520
rect 121656 700262 121684 703520
rect 137848 702434 137876 703520
rect 137848 702406 137968 702434
rect 121644 700256 121696 700262
rect 121644 700198 121696 700204
rect 122748 700256 122800 700262
rect 122748 700198 122800 700204
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 99288 369368 99340 369374
rect 99288 369310 99340 369316
rect 89628 369232 89680 369238
rect 89628 369174 89680 369180
rect 99300 366194 99328 369310
rect 106200 369306 106228 699654
rect 106188 369300 106240 369306
rect 106188 369242 106240 369248
rect 118976 369232 119028 369238
rect 118976 369174 119028 369180
rect 109132 369164 109184 369170
rect 109132 369106 109184 369112
rect 109144 366194 109172 369106
rect 118988 366194 119016 369174
rect 122760 369170 122788 700198
rect 128820 369300 128872 369306
rect 128820 369242 128872 369248
rect 122748 369164 122800 369170
rect 122748 369106 122800 369112
rect 128832 366194 128860 369242
rect 137940 369238 137968 702406
rect 154132 700126 154160 703520
rect 154120 700120 154172 700126
rect 154120 700062 154172 700068
rect 155224 700120 155276 700126
rect 155224 700062 155276 700068
rect 155236 369238 155264 700062
rect 170324 699718 170352 703520
rect 186516 700398 186544 703520
rect 202800 700466 202828 703520
rect 217968 700596 218020 700602
rect 217968 700538 218020 700544
rect 188988 700460 189040 700466
rect 188988 700402 189040 700408
rect 202788 700460 202840 700466
rect 202788 700402 202840 700408
rect 177948 700392 178000 700398
rect 177948 700334 178000 700340
rect 186504 700392 186556 700398
rect 186504 700334 186556 700340
rect 169024 699712 169076 699718
rect 169024 699654 169076 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 169036 369850 169064 699654
rect 168104 369844 168156 369850
rect 168104 369786 168156 369792
rect 169024 369844 169076 369850
rect 169024 369786 169076 369792
rect 137928 369232 137980 369238
rect 137928 369174 137980 369180
rect 148416 369232 148468 369238
rect 148416 369174 148468 369180
rect 155224 369232 155276 369238
rect 155224 369174 155276 369180
rect 158260 369232 158312 369238
rect 158260 369174 158312 369180
rect 138572 369164 138624 369170
rect 138572 369106 138624 369112
rect 60844 366166 60888 366194
rect 69768 366166 69845 366194
rect 79612 366166 79676 366194
rect 89456 366166 89506 366194
rect 99300 366166 99337 366194
rect 60860 365915 60888 366166
rect 69817 365915 69845 366166
rect 79648 365915 79676 366166
rect 89478 365915 89506 366166
rect 99309 365915 99337 366166
rect 109140 366166 109172 366194
rect 118971 366166 119016 366194
rect 128802 366166 128860 366194
rect 109140 365915 109168 366166
rect 118971 365915 118999 366166
rect 128802 365915 128830 366166
rect 138584 366058 138612 369106
rect 148428 366194 148456 369174
rect 158272 366194 158300 369174
rect 168116 366194 168144 369786
rect 177960 366194 177988 700334
rect 189000 369170 189028 700402
rect 198648 700392 198700 700398
rect 198648 700334 198700 700340
rect 198660 369714 198688 700334
rect 217980 369850 218008 700538
rect 218992 700398 219020 703520
rect 227628 700528 227680 700534
rect 227628 700470 227680 700476
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 220084 700392 220136 700398
rect 220084 700334 220136 700340
rect 217232 369844 217284 369850
rect 217232 369786 217284 369792
rect 217968 369844 218020 369850
rect 217968 369786 218020 369792
rect 197636 369708 197688 369714
rect 197636 369650 197688 369656
rect 198648 369708 198700 369714
rect 198648 369650 198700 369656
rect 187792 369164 187844 369170
rect 187792 369106 187844 369112
rect 188988 369164 189040 369170
rect 188988 369106 189040 369112
rect 187804 366194 187832 369106
rect 197648 366194 197676 369650
rect 207480 369164 207532 369170
rect 207480 369106 207532 369112
rect 148428 366166 148491 366194
rect 158272 366166 158322 366194
rect 168116 366166 168153 366194
rect 138584 366030 138660 366058
rect 138632 365915 138660 366030
rect 148463 365915 148491 366166
rect 158294 365915 158322 366166
rect 168125 365915 168153 366166
rect 177956 366166 177988 366194
rect 187786 366166 187832 366194
rect 197617 366166 197676 366194
rect 177956 365915 177984 366166
rect 187786 365915 187814 366166
rect 197617 365915 197645 366166
rect 207492 366058 207520 369106
rect 217244 366194 217272 369786
rect 220096 369170 220124 700334
rect 227640 369850 227668 700470
rect 235184 700398 235212 703520
rect 251468 700602 251496 703520
rect 256608 700732 256660 700738
rect 256608 700674 256660 700680
rect 251456 700596 251508 700602
rect 251456 700538 251508 700544
rect 237288 700460 237340 700466
rect 237288 700402 237340 700408
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 237300 373994 237328 700402
rect 246948 700392 247000 700398
rect 246948 700334 247000 700340
rect 246960 373994 246988 700334
rect 237024 373966 237328 373994
rect 246776 373966 246988 373994
rect 227076 369844 227128 369850
rect 227076 369786 227128 369792
rect 227628 369844 227680 369850
rect 227628 369786 227680 369792
rect 220084 369164 220136 369170
rect 220084 369106 220136 369112
rect 227088 366194 227116 369786
rect 237024 366194 237052 373966
rect 246776 366194 246804 373966
rect 256620 366194 256648 700674
rect 267556 700664 267608 700670
rect 267556 700606 267608 700612
rect 267568 692774 267596 700606
rect 267660 700534 267688 703520
rect 277308 700596 277360 700602
rect 277308 700538 277360 700544
rect 267648 700528 267700 700534
rect 267648 700470 267700 700476
rect 267568 692746 267688 692774
rect 267660 369102 267688 692746
rect 266452 369096 266504 369102
rect 266452 369038 266504 369044
rect 267648 369096 267700 369102
rect 267648 369038 267700 369044
rect 266464 366194 266492 369038
rect 277320 369034 277348 700538
rect 283852 700466 283880 703520
rect 286968 700528 287020 700534
rect 286968 700470 287020 700476
rect 283840 700460 283892 700466
rect 283840 700402 283892 700408
rect 286980 369850 287008 700470
rect 296628 700460 296680 700466
rect 296628 700402 296680 700408
rect 296640 369850 296668 700402
rect 300136 700398 300164 703520
rect 315948 701004 316000 701010
rect 315948 700946 316000 700952
rect 300124 700392 300176 700398
rect 300124 700334 300176 700340
rect 306288 700392 306340 700398
rect 306288 700334 306340 700340
rect 306300 369850 306328 700334
rect 315960 373994 315988 700946
rect 316328 700738 316356 703520
rect 325608 700936 325660 700942
rect 325608 700878 325660 700884
rect 316316 700732 316368 700738
rect 316316 700674 316368 700680
rect 325620 373994 325648 700878
rect 332520 700670 332548 703520
rect 335268 700868 335320 700874
rect 335268 700810 335320 700816
rect 332508 700664 332560 700670
rect 332508 700606 332560 700612
rect 315592 373966 315988 373994
rect 325436 373966 325648 373994
rect 286048 369844 286100 369850
rect 286048 369786 286100 369792
rect 286968 369844 287020 369850
rect 286968 369786 287020 369792
rect 295892 369844 295944 369850
rect 295892 369786 295944 369792
rect 296628 369844 296680 369850
rect 296628 369786 296680 369792
rect 305736 369844 305788 369850
rect 305736 369786 305788 369792
rect 306288 369844 306340 369850
rect 306288 369786 306340 369792
rect 276296 369028 276348 369034
rect 276296 368970 276348 368976
rect 277308 369028 277360 369034
rect 277308 368970 277360 368976
rect 217244 366166 217307 366194
rect 227088 366166 227138 366194
rect 207448 366030 207520 366058
rect 207448 365915 207476 366030
rect 217279 365915 217307 366166
rect 227110 365915 227138 366166
rect 236940 366166 237052 366194
rect 246771 366166 246804 366194
rect 256602 366166 256648 366194
rect 266433 366166 266492 366194
rect 236940 365915 236968 366166
rect 246771 365915 246799 366166
rect 256602 365915 256630 366166
rect 266433 365915 266461 366166
rect 276308 366058 276336 368970
rect 286060 366194 286088 369786
rect 295904 366194 295932 369786
rect 305748 366194 305776 369786
rect 315592 366194 315620 373966
rect 325436 366194 325464 373966
rect 335280 366194 335308 700810
rect 346308 700800 346360 700806
rect 346308 700742 346360 700748
rect 346320 369170 346348 700742
rect 348804 700602 348832 703520
rect 355968 700732 356020 700738
rect 355968 700674 356020 700680
rect 348792 700596 348844 700602
rect 348792 700538 348844 700544
rect 355980 369850 356008 700674
rect 364996 700534 365024 703520
rect 365628 700664 365680 700670
rect 365628 700606 365680 700612
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 365640 369850 365668 700606
rect 375288 700596 375340 700602
rect 375288 700538 375340 700544
rect 375300 369850 375328 700538
rect 381188 700466 381216 703520
rect 384948 700528 385000 700534
rect 384948 700470 385000 700476
rect 381176 700460 381228 700466
rect 381176 700402 381228 700408
rect 384960 369850 384988 700470
rect 394608 700460 394660 700466
rect 394608 700402 394660 700408
rect 394620 373994 394648 700402
rect 397472 700398 397500 703520
rect 413664 701010 413692 703520
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 429856 700942 429884 703520
rect 429844 700936 429896 700942
rect 429844 700878 429896 700884
rect 446140 700874 446168 703520
rect 446128 700868 446180 700874
rect 446128 700810 446180 700816
rect 462332 700806 462360 703520
rect 462320 700800 462372 700806
rect 462320 700742 462372 700748
rect 478524 700738 478552 703520
rect 478512 700732 478564 700738
rect 478512 700674 478564 700680
rect 494808 700670 494836 703520
rect 494796 700664 494848 700670
rect 494796 700606 494848 700612
rect 511000 700602 511028 703520
rect 510988 700596 511040 700602
rect 510988 700538 511040 700544
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 700398 559696 703520
rect 397460 700392 397512 700398
rect 397460 700334 397512 700340
rect 404268 700392 404320 700398
rect 404268 700334 404320 700340
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 394252 373966 394648 373994
rect 354864 369844 354916 369850
rect 354864 369786 354916 369792
rect 355968 369844 356020 369850
rect 355968 369786 356020 369792
rect 364708 369844 364760 369850
rect 364708 369786 364760 369792
rect 365628 369844 365680 369850
rect 365628 369786 365680 369792
rect 374552 369844 374604 369850
rect 374552 369786 374604 369792
rect 375288 369844 375340 369850
rect 375288 369786 375340 369792
rect 384396 369844 384448 369850
rect 384396 369786 384448 369792
rect 384948 369844 385000 369850
rect 384948 369786 385000 369792
rect 345112 369164 345164 369170
rect 345112 369106 345164 369112
rect 346308 369164 346360 369170
rect 346308 369106 346360 369112
rect 286060 366166 286122 366194
rect 295904 366166 295953 366194
rect 305748 366166 305784 366194
rect 276264 366030 276336 366058
rect 276264 365915 276292 366030
rect 286094 365915 286122 366166
rect 295925 365915 295953 366166
rect 305756 365915 305784 366166
rect 315587 366166 315620 366194
rect 325418 366166 325464 366194
rect 335248 366166 335308 366194
rect 315587 365915 315615 366166
rect 325418 365915 325446 366166
rect 335248 365915 335276 366166
rect 345124 366058 345152 369106
rect 354876 366194 354904 369786
rect 364720 366194 364748 369786
rect 374564 366194 374592 369786
rect 384408 366194 384436 369786
rect 394252 366194 394280 373966
rect 404280 369850 404308 700334
rect 575860 700330 575888 703520
rect 575848 700324 575900 700330
rect 575848 700266 575900 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 411904 696992 411956 696998
rect 411904 696934 411956 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 406384 683188 406436 683194
rect 406384 683130 406436 683136
rect 406292 418192 406344 418198
rect 406292 418134 406344 418140
rect 406200 404388 406252 404394
rect 406200 404330 406252 404336
rect 406108 378208 406160 378214
rect 406108 378150 406160 378156
rect 402980 369844 403032 369850
rect 402980 369786 403032 369792
rect 404268 369844 404320 369850
rect 404268 369786 404320 369792
rect 354876 366166 354938 366194
rect 364720 366166 364769 366194
rect 374564 366166 374600 366194
rect 345079 366030 345152 366058
rect 345079 365915 345107 366030
rect 354910 365915 354938 366166
rect 364741 365915 364769 366166
rect 374572 365915 374600 366166
rect 384402 366166 384436 366194
rect 394233 366166 394280 366194
rect 402992 366194 403020 369786
rect 402992 366166 403036 366194
rect 384402 365915 384430 366166
rect 394233 365915 394261 366166
rect 403008 365915 403036 366166
rect 57428 365696 57480 365702
rect 57428 365638 57480 365644
rect 57440 365129 57468 365638
rect 57426 365120 57482 365129
rect 57426 365055 57482 365064
rect 406016 365016 406068 365022
rect 406014 364984 406016 364993
rect 406068 364984 406070 364993
rect 406014 364919 406070 364928
rect 57152 361548 57204 361554
rect 57152 361490 57204 361496
rect 57164 360505 57192 361490
rect 57150 360496 57206 360505
rect 57150 360431 57206 360440
rect 57244 356040 57296 356046
rect 57244 355982 57296 355988
rect 57256 354929 57284 355982
rect 57242 354920 57298 354929
rect 57242 354855 57298 354864
rect 57612 350532 57664 350538
rect 57612 350474 57664 350480
rect 57624 349353 57652 350474
rect 57610 349344 57666 349353
rect 57610 349279 57666 349288
rect 57612 345024 57664 345030
rect 57612 344966 57664 344972
rect 57624 343777 57652 344966
rect 57610 343768 57666 343777
rect 57610 343703 57666 343712
rect 57612 339448 57664 339454
rect 57612 339390 57664 339396
rect 57624 338337 57652 339390
rect 57610 338328 57666 338337
rect 57610 338263 57666 338272
rect 57612 333940 57664 333946
rect 57612 333882 57664 333888
rect 57624 332761 57652 333882
rect 57610 332752 57666 332761
rect 57610 332687 57666 332696
rect 57336 328432 57388 328438
rect 57336 328374 57388 328380
rect 57348 327185 57376 328374
rect 57334 327176 57390 327185
rect 57334 327111 57390 327120
rect 57336 322924 57388 322930
rect 57336 322866 57388 322872
rect 57348 321609 57376 322866
rect 57334 321600 57390 321609
rect 57334 321535 57390 321544
rect 57612 317416 57664 317422
rect 57612 317358 57664 317364
rect 57624 316169 57652 317358
rect 57610 316160 57666 316169
rect 57610 316095 57666 316104
rect 57612 310480 57664 310486
rect 57610 310448 57612 310457
rect 57664 310448 57666 310457
rect 57610 310383 57666 310392
rect 57426 305008 57482 305017
rect 57426 304943 57428 304952
rect 57480 304943 57482 304952
rect 57428 304914 57480 304920
rect 57612 299464 57664 299470
rect 57610 299432 57612 299441
rect 57664 299432 57666 299441
rect 57610 299367 57666 299376
rect 405832 299328 405884 299334
rect 405832 299270 405884 299276
rect 405844 298217 405872 299270
rect 405830 298208 405886 298217
rect 405830 298143 405886 298152
rect 57612 293956 57664 293962
rect 57612 293898 57664 293904
rect 57624 293865 57652 293898
rect 57610 293856 57666 293865
rect 57610 293791 57666 293800
rect 57610 288416 57666 288425
rect 57610 288351 57612 288360
rect 57664 288351 57666 288360
rect 57612 288322 57664 288328
rect 57612 282872 57664 282878
rect 57610 282840 57612 282849
rect 57664 282840 57666 282849
rect 57610 282775 57666 282784
rect 57612 277364 57664 277370
rect 57612 277306 57664 277312
rect 57624 277273 57652 277306
rect 57610 277264 57666 277273
rect 57610 277199 57666 277208
rect 57520 271856 57572 271862
rect 57520 271798 57572 271804
rect 57532 271697 57560 271798
rect 57518 271688 57574 271697
rect 57518 271623 57574 271632
rect 39304 266348 39356 266354
rect 39304 266290 39356 266296
rect 57336 266348 57388 266354
rect 57336 266290 57388 266296
rect 57348 266121 57376 266290
rect 57334 266112 57390 266121
rect 57334 266047 57390 266056
rect 33784 260840 33836 260846
rect 33784 260782 33836 260788
rect 57428 260840 57480 260846
rect 57428 260782 57480 260788
rect 57440 260681 57468 260782
rect 57426 260672 57482 260681
rect 57426 260607 57482 260616
rect 57612 255264 57664 255270
rect 57612 255206 57664 255212
rect 57624 255105 57652 255206
rect 57610 255096 57666 255105
rect 57610 255031 57666 255040
rect 21364 249756 21416 249762
rect 21364 249698 21416 249704
rect 57244 249756 57296 249762
rect 57244 249698 57296 249704
rect 57256 249529 57284 249698
rect 57242 249520 57298 249529
rect 57242 249455 57298 249464
rect 57428 244248 57480 244254
rect 57428 244190 57480 244196
rect 57440 243953 57468 244190
rect 57426 243944 57482 243953
rect 57426 243879 57482 243888
rect 4068 238740 4120 238746
rect 4068 238682 4120 238688
rect 57612 238740 57664 238746
rect 57612 238682 57664 238688
rect 57624 238513 57652 238682
rect 57610 238504 57666 238513
rect 57610 238439 57666 238448
rect 57612 233232 57664 233238
rect 57612 233174 57664 233180
rect 57624 232937 57652 233174
rect 57610 232928 57666 232937
rect 57610 232863 57666 232872
rect 406120 230353 406148 378150
rect 406212 241641 406240 404330
rect 406304 247217 406332 418134
rect 406396 360369 406424 683130
rect 406476 670744 406528 670750
rect 406476 670686 406528 670692
rect 406382 360360 406438 360369
rect 406382 360295 406438 360304
rect 406488 354657 406516 670686
rect 410524 643136 410576 643142
rect 410524 643078 410576 643084
rect 406568 616888 406620 616894
rect 406568 616830 406620 616836
rect 406474 354648 406530 354657
rect 406474 354583 406530 354592
rect 406384 351960 406436 351966
rect 406384 351902 406436 351908
rect 406290 247208 406346 247217
rect 406290 247143 406346 247152
rect 406198 241632 406254 241641
rect 406198 241567 406254 241576
rect 406106 230344 406162 230353
rect 406106 230279 406162 230288
rect 3974 228032 4030 228041
rect 3974 227967 4030 227976
rect 3884 172508 3936 172514
rect 3884 172450 3936 172456
rect 3988 167006 4016 227967
rect 57612 227724 57664 227730
rect 57612 227666 57664 227672
rect 57624 227361 57652 227666
rect 57610 227352 57666 227361
rect 57610 227287 57666 227296
rect 406292 224664 406344 224670
rect 406290 224632 406292 224641
rect 406344 224632 406346 224641
rect 406290 224567 406346 224576
rect 57612 222148 57664 222154
rect 57612 222090 57664 222096
rect 57624 221785 57652 222090
rect 57610 221776 57666 221785
rect 57610 221711 57666 221720
rect 406396 219065 406424 351902
rect 406476 349104 406528 349110
rect 406474 349072 406476 349081
rect 406528 349072 406530 349081
rect 406474 349007 406530 349016
rect 406476 343392 406528 343398
rect 406474 343360 406476 343369
rect 406528 343360 406530 343369
rect 406474 343295 406530 343304
rect 406476 338088 406528 338094
rect 406476 338030 406528 338036
rect 406488 337793 406516 338030
rect 406474 337784 406530 337793
rect 406474 337719 406530 337728
rect 406580 335354 406608 616830
rect 406660 590708 406712 590714
rect 406660 590650 406712 590656
rect 406488 335326 406608 335354
rect 406488 332081 406516 335326
rect 406474 332072 406530 332081
rect 406474 332007 406530 332016
rect 406568 327072 406620 327078
rect 406568 327014 406620 327020
rect 406580 326369 406608 327014
rect 406566 326360 406622 326369
rect 406566 326295 406622 326304
rect 406476 324352 406528 324358
rect 406476 324294 406528 324300
rect 406382 219056 406438 219065
rect 406382 218991 406438 219000
rect 406292 218068 406344 218074
rect 406292 218010 406344 218016
rect 57060 216640 57112 216646
rect 57060 216582 57112 216588
rect 57072 216209 57100 216582
rect 57058 216200 57114 216209
rect 57058 216135 57114 216144
rect 56784 211132 56836 211138
rect 56784 211074 56836 211080
rect 56796 210769 56824 211074
rect 56782 210760 56838 210769
rect 56782 210695 56838 210704
rect 57612 205624 57664 205630
rect 57612 205566 57664 205572
rect 57624 205193 57652 205566
rect 57610 205184 57666 205193
rect 57610 205119 57666 205128
rect 57612 200116 57664 200122
rect 57612 200058 57664 200064
rect 57624 199617 57652 200058
rect 57610 199608 57666 199617
rect 57610 199543 57666 199552
rect 57612 194540 57664 194546
rect 57612 194482 57664 194488
rect 57624 194041 57652 194482
rect 57610 194032 57666 194041
rect 57610 193967 57666 193976
rect 57612 189032 57664 189038
rect 57612 188974 57664 188980
rect 57624 188601 57652 188974
rect 57610 188592 57666 188601
rect 57610 188527 57666 188536
rect 57612 183524 57664 183530
rect 57612 183466 57664 183472
rect 57624 183025 57652 183466
rect 57610 183016 57666 183025
rect 57610 182951 57666 182960
rect 56692 178016 56744 178022
rect 56692 177958 56744 177964
rect 56704 177449 56732 177958
rect 56690 177440 56746 177449
rect 56690 177375 56746 177384
rect 57612 172508 57664 172514
rect 57612 172450 57664 172456
rect 57624 171873 57652 172450
rect 57610 171864 57666 171873
rect 57610 171799 57666 171808
rect 3976 167000 4028 167006
rect 3976 166942 4028 166948
rect 57612 167000 57664 167006
rect 57612 166942 57664 166948
rect 57624 166297 57652 166942
rect 57610 166288 57666 166297
rect 57610 166223 57666 166232
rect 3790 162888 3846 162897
rect 3790 162823 3846 162832
rect 3700 144900 3752 144906
rect 3700 144842 3752 144848
rect 3804 139398 3832 162823
rect 406304 162489 406332 218010
rect 406384 213920 406436 213926
rect 406384 213862 406436 213868
rect 406396 213353 406424 213862
rect 406382 213344 406438 213353
rect 406382 213279 406438 213288
rect 406488 207777 406516 324294
rect 406672 320793 406700 590650
rect 406752 576904 406804 576910
rect 406752 576846 406804 576852
rect 406658 320784 406714 320793
rect 406658 320719 406714 320728
rect 406764 315081 406792 576846
rect 406844 563100 406896 563106
rect 406844 563042 406896 563048
rect 406750 315072 406806 315081
rect 406750 315007 406806 315016
rect 406568 311908 406620 311914
rect 406568 311850 406620 311856
rect 406474 207768 406530 207777
rect 406474 207703 406530 207712
rect 406384 205692 406436 205698
rect 406384 205634 406436 205640
rect 406290 162480 406346 162489
rect 406290 162415 406346 162424
rect 57612 161424 57664 161430
rect 57612 161366 57664 161372
rect 57624 160857 57652 161366
rect 57610 160848 57666 160857
rect 57610 160783 57666 160792
rect 406396 156777 406424 205634
rect 406580 202065 406608 311850
rect 406856 309505 406884 563042
rect 407764 536852 407816 536858
rect 407764 536794 407816 536800
rect 406936 484424 406988 484430
rect 406936 484366 406988 484372
rect 406842 309496 406898 309505
rect 406842 309431 406898 309440
rect 406844 304972 406896 304978
rect 406844 304914 406896 304920
rect 406856 303793 406884 304914
rect 406842 303784 406898 303793
rect 406842 303719 406898 303728
rect 406660 298172 406712 298178
rect 406660 298114 406712 298120
rect 406566 202056 406622 202065
rect 406566 201991 406622 202000
rect 406672 196353 406700 298114
rect 406844 292528 406896 292534
rect 406842 292496 406844 292505
rect 406896 292496 406898 292505
rect 406842 292431 406898 292440
rect 406844 287020 406896 287026
rect 406844 286962 406896 286968
rect 406856 286793 406884 286962
rect 406842 286784 406898 286793
rect 406842 286719 406898 286728
rect 406844 281512 406896 281518
rect 406844 281454 406896 281460
rect 406856 281217 406884 281454
rect 406842 281208 406898 281217
rect 406842 281143 406898 281152
rect 406948 275505 406976 484366
rect 407028 470620 407080 470626
rect 407028 470562 407080 470568
rect 406934 275496 406990 275505
rect 406934 275431 406990 275440
rect 406752 271924 406804 271930
rect 406752 271866 406804 271872
rect 406658 196344 406714 196353
rect 406658 196279 406714 196288
rect 406764 195242 406792 271866
rect 407040 269929 407068 470562
rect 407776 299334 407804 536794
rect 410536 343398 410564 643078
rect 411916 365022 411944 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580262 657384 580318 657393
rect 580262 657319 580318 657328
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 418804 630692 418856 630698
rect 418804 630634 418856 630640
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 417424 524476 417476 524482
rect 417424 524418 417476 524424
rect 414664 430636 414716 430642
rect 414664 430578 414716 430584
rect 411904 365016 411956 365022
rect 411904 364958 411956 364964
rect 411996 364404 412048 364410
rect 411996 364346 412048 364352
rect 410524 343392 410576 343398
rect 410524 343334 410576 343340
rect 407764 299328 407816 299334
rect 407764 299270 407816 299276
rect 407026 269920 407082 269929
rect 407026 269855 407082 269864
rect 407028 264920 407080 264926
rect 407028 264862 407080 264868
rect 407040 264217 407068 264862
rect 407026 264208 407082 264217
rect 407026 264143 407082 264152
rect 406936 259412 406988 259418
rect 406936 259354 406988 259360
rect 406844 258120 406896 258126
rect 406948 258097 406976 259354
rect 406844 258062 406896 258068
rect 406934 258088 406990 258097
rect 406672 195214 406792 195242
rect 406476 191888 406528 191894
rect 406476 191830 406528 191836
rect 406382 156768 406438 156777
rect 406382 156703 406438 156712
rect 57612 155916 57664 155922
rect 57612 155858 57664 155864
rect 57624 155281 57652 155858
rect 57610 155272 57666 155281
rect 57610 155207 57666 155216
rect 406384 151836 406436 151842
rect 406384 151778 406436 151784
rect 56876 150408 56928 150414
rect 56876 150350 56928 150356
rect 56888 149705 56916 150350
rect 56874 149696 56930 149705
rect 56874 149631 56930 149640
rect 57520 144900 57572 144906
rect 57520 144842 57572 144848
rect 57532 144129 57560 144842
rect 57518 144120 57574 144129
rect 57518 144055 57574 144064
rect 3792 139392 3844 139398
rect 3792 139334 3844 139340
rect 57520 139392 57572 139398
rect 57520 139334 57572 139340
rect 57532 138553 57560 139334
rect 57518 138544 57574 138553
rect 57518 138479 57574 138488
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3424 133884 3476 133890
rect 3424 133826 3476 133832
rect 3528 128314 3556 136711
rect 406396 134201 406424 151778
rect 406488 151201 406516 191830
rect 406672 185065 406700 195214
rect 406752 191820 406804 191826
rect 406752 191762 406804 191768
rect 406764 190777 406792 191762
rect 406750 190768 406806 190777
rect 406750 190703 406806 190712
rect 406658 185056 406714 185065
rect 406658 184991 406714 185000
rect 406856 179489 406884 258062
rect 406934 258023 406990 258032
rect 407026 252920 407082 252929
rect 407026 252855 407028 252864
rect 407080 252855 407082 252864
rect 407028 252826 407080 252832
rect 406936 244316 406988 244322
rect 406936 244258 406988 244264
rect 406842 179480 406898 179489
rect 406842 179415 406898 179424
rect 406568 178084 406620 178090
rect 406568 178026 406620 178032
rect 406474 151192 406530 151201
rect 406474 151127 406530 151136
rect 406580 145489 406608 178026
rect 406948 173777 406976 244258
rect 407028 235952 407080 235958
rect 407026 235920 407028 235929
rect 407080 235920 407082 235929
rect 407026 235855 407082 235864
rect 407028 231872 407080 231878
rect 407028 231814 407080 231820
rect 406934 173768 406990 173777
rect 406934 173703 406990 173712
rect 407040 168201 407068 231814
rect 412008 224670 412036 364346
rect 414676 252890 414704 430578
rect 417436 292534 417464 524418
rect 418816 338094 418844 630634
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579618 591016 579674 591025
rect 579618 590951 579674 590960
rect 579632 590714 579660 590951
rect 579620 590708 579672 590714
rect 579620 590650 579672 590656
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 576910 579660 577623
rect 579620 576904 579672 576910
rect 579620 576846 579672 576852
rect 579894 564360 579950 564369
rect 579894 564295 579950 564304
rect 579908 563106 579936 564295
rect 579896 563100 579948 563106
rect 579896 563042 579948 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 579618 484664 579674 484673
rect 579618 484599 579674 484608
rect 579632 484430 579660 484599
rect 579620 484424 579672 484430
rect 579620 484366 579672 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 579986 431624 580042 431633
rect 579986 431559 580042 431568
rect 580000 430642 580028 431559
rect 579988 430636 580040 430642
rect 579988 430578 580040 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 579816 378214 579844 378383
rect 579804 378208 579856 378214
rect 579804 378150 579856 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580276 354674 580304 657319
rect 580354 604208 580410 604217
rect 580354 604143 580410 604152
rect 580092 354646 580304 354674
rect 580092 349110 580120 354646
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580080 349104 580132 349110
rect 580080 349046 580132 349052
rect 580262 338600 580318 338609
rect 580262 338535 580318 338544
rect 418804 338088 418856 338094
rect 418804 338030 418856 338036
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 417424 292528 417476 292534
rect 417424 292470 417476 292476
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 414664 252884 414716 252890
rect 414664 252826 414716 252832
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 579632 231878 579660 232319
rect 579620 231872 579672 231878
rect 579620 231814 579672 231820
rect 411996 224664 412048 224670
rect 411996 224606 412048 224612
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 580276 213926 580304 338535
rect 580368 327078 580396 604143
rect 580446 551168 580502 551177
rect 580446 551103 580502 551112
rect 580356 327072 580408 327078
rect 580356 327014 580408 327020
rect 580460 304978 580488 551103
rect 580538 511320 580594 511329
rect 580538 511255 580594 511264
rect 580448 304972 580500 304978
rect 580448 304914 580500 304920
rect 580552 287026 580580 511255
rect 580630 497992 580686 498001
rect 580630 497927 580686 497936
rect 580540 287020 580592 287026
rect 580540 286962 580592 286968
rect 580354 285424 580410 285433
rect 580354 285359 580410 285368
rect 580264 213920 580316 213926
rect 580264 213862 580316 213868
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 580368 191826 580396 285359
rect 580644 281518 580672 497927
rect 580722 458144 580778 458153
rect 580722 458079 580778 458088
rect 580632 281512 580684 281518
rect 580632 281454 580684 281460
rect 580736 264926 580764 458079
rect 580814 444816 580870 444825
rect 580814 444751 580870 444760
rect 580724 264920 580776 264926
rect 580724 264862 580776 264868
rect 580828 259418 580856 444751
rect 580906 391776 580962 391785
rect 580906 391711 580962 391720
rect 580816 259412 580868 259418
rect 580816 259354 580868 259360
rect 580920 235958 580948 391711
rect 580908 235952 580960 235958
rect 580908 235894 580960 235900
rect 580356 191820 580408 191826
rect 580356 191762 580408 191768
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 407026 168192 407082 168201
rect 407026 168127 407082 168136
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 406660 165640 406712 165646
rect 406660 165582 406712 165588
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 406566 145480 406622 145489
rect 406566 145415 406622 145424
rect 406672 139913 406700 165582
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 406658 139904 406714 139913
rect 406658 139839 406714 139848
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 406476 138032 406528 138038
rect 406476 137974 406528 137980
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 406382 134192 406438 134201
rect 406382 134127 406438 134136
rect 57520 133884 57572 133890
rect 57520 133826 57572 133832
rect 57532 133113 57560 133826
rect 57518 133104 57574 133113
rect 57518 133039 57574 133048
rect 406488 128625 406516 137974
rect 406474 128616 406530 128625
rect 406474 128551 406530 128560
rect 3516 128308 3568 128314
rect 3516 128250 3568 128256
rect 56968 128308 57020 128314
rect 56968 128250 57020 128256
rect 56980 127537 57008 128250
rect 56966 127528 57022 127537
rect 56966 127463 57022 127472
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580184 125662 580212 125967
rect 407028 125656 407080 125662
rect 407028 125598 407080 125604
rect 580172 125656 580224 125662
rect 580172 125598 580224 125604
rect 3606 123720 3662 123729
rect 3606 123655 3662 123664
rect 3620 122806 3648 123655
rect 407040 122913 407068 125598
rect 407026 122904 407082 122913
rect 407026 122839 407082 122848
rect 3608 122800 3660 122806
rect 3608 122742 3660 122748
rect 57060 122800 57112 122806
rect 57060 122742 57112 122748
rect 57072 121961 57100 122742
rect 57058 121952 57114 121961
rect 57058 121887 57114 121896
rect 406382 117192 406438 117201
rect 406382 117127 406438 117136
rect 57610 116376 57666 116385
rect 57610 116311 57666 116320
rect 57624 116006 57652 116311
rect 3424 116000 3476 116006
rect 3424 115942 3476 115948
rect 57612 116000 57664 116006
rect 57612 115942 57664 115948
rect 3436 110673 3464 115942
rect 406396 113150 406424 117127
rect 406384 113144 406436 113150
rect 406384 113086 406436 113092
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 406474 111616 406530 111625
rect 406474 111551 406530 111560
rect 57610 110800 57666 110809
rect 57610 110735 57666 110744
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 57624 110498 57652 110735
rect 3516 110492 3568 110498
rect 3516 110434 3568 110440
rect 57612 110492 57664 110498
rect 57612 110434 57664 110440
rect 3424 104916 3476 104922
rect 3424 104858 3476 104864
rect 3436 84697 3464 104858
rect 3528 97617 3556 110434
rect 406382 105904 406438 105913
rect 406382 105839 406438 105848
rect 57426 105224 57482 105233
rect 57426 105159 57482 105168
rect 57440 104922 57468 105159
rect 57428 104916 57480 104922
rect 57428 104858 57480 104864
rect 57426 99784 57482 99793
rect 57426 99719 57482 99728
rect 57440 99414 57468 99719
rect 3884 99408 3936 99414
rect 3884 99350 3936 99356
rect 57428 99408 57480 99414
rect 57428 99350 57480 99356
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3792 93900 3844 93906
rect 3792 93842 3844 93848
rect 3700 88392 3752 88398
rect 3700 88334 3752 88340
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3608 82884 3660 82890
rect 3608 82826 3660 82832
rect 3516 77308 3568 77314
rect 3516 77250 3568 77256
rect 3424 71800 3476 71806
rect 3424 71742 3476 71748
rect 3436 6497 3464 71742
rect 3528 19417 3556 77250
rect 3620 32473 3648 82826
rect 3712 45529 3740 88334
rect 3804 58585 3832 93842
rect 3896 71641 3924 99350
rect 57610 94208 57666 94217
rect 57610 94143 57666 94152
rect 57624 93906 57652 94143
rect 57612 93900 57664 93906
rect 57612 93842 57664 93848
rect 57518 88632 57574 88641
rect 57518 88567 57574 88576
rect 57532 88398 57560 88567
rect 57520 88392 57572 88398
rect 57520 88334 57572 88340
rect 406396 86970 406424 105839
rect 406488 100706 406516 111551
rect 406476 100700 406528 100706
rect 406476 100642 406528 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 406842 100328 406898 100337
rect 406842 100263 406898 100272
rect 406750 94616 406806 94625
rect 406750 94551 406806 94560
rect 406658 88904 406714 88913
rect 406658 88839 406714 88848
rect 406384 86964 406436 86970
rect 406384 86906 406436 86912
rect 406566 83328 406622 83337
rect 406566 83263 406622 83272
rect 57426 83056 57482 83065
rect 57426 82991 57482 83000
rect 57440 82890 57468 82991
rect 57428 82884 57480 82890
rect 57428 82826 57480 82832
rect 57518 77616 57574 77625
rect 57518 77551 57574 77560
rect 406474 77616 406530 77625
rect 406474 77551 406530 77560
rect 57532 77314 57560 77551
rect 57520 77308 57572 77314
rect 57520 77250 57572 77256
rect 57426 72856 57482 72865
rect 57426 72791 57482 72800
rect 406382 72856 406438 72865
rect 406382 72791 406438 72800
rect 57440 71806 57468 72791
rect 57428 71800 57480 71806
rect 60308 71754 60336 72012
rect 60684 71754 60712 72012
rect 57428 71742 57480 71748
rect 60292 71726 60336 71754
rect 60660 71726 60712 71754
rect 60832 71800 60884 71806
rect 60832 71742 60884 71748
rect 61382 71754 61410 72012
rect 62079 71806 62107 72012
rect 62067 71800 62119 71806
rect 3882 71632 3938 71641
rect 3882 71567 3938 71576
rect 53104 70372 53156 70378
rect 53104 70314 53156 70320
rect 41328 70304 41380 70310
rect 41328 70246 41380 70252
rect 34428 70236 34480 70242
rect 34428 70178 34480 70184
rect 27528 70100 27580 70106
rect 27528 70042 27580 70048
rect 17868 69964 17920 69970
rect 17868 69906 17920 69912
rect 7564 69896 7616 69902
rect 7564 69838 7616 69844
rect 3790 58576 3846 58585
rect 3790 58511 3846 58520
rect 3698 45520 3754 45529
rect 3698 45455 3754 45464
rect 3606 32464 3662 32473
rect 3606 32399 3662 32408
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 6190
rect 4068 4956 4120 4962
rect 4068 4898 4120 4904
rect 4080 480 4108 4898
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 3538
rect 7576 3466 7604 69838
rect 11704 69692 11756 69698
rect 11704 69634 11756 69640
rect 7656 4888 7708 4894
rect 7656 4830 7708 4836
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7668 480 7696 4830
rect 11716 3602 11744 69634
rect 14464 68604 14516 68610
rect 14464 68546 14516 68552
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 11150 3496 11206 3505
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8772 480 8800 3402
rect 9968 480 9996 3470
rect 11150 3431 11206 3440
rect 11164 480 11192 3431
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12360 480 12388 3062
rect 13556 480 13584 3538
rect 14476 3126 14504 68546
rect 15844 66904 15896 66910
rect 15844 66846 15896 66852
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14752 480 14780 3946
rect 15856 3534 15884 66846
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15948 480 15976 3606
rect 17880 3534 17908 69906
rect 18604 69828 18656 69834
rect 18604 69770 18656 69776
rect 18616 4010 18644 69770
rect 21364 69760 21416 69766
rect 21364 69702 21416 69708
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 21376 3670 21404 69702
rect 25504 68468 25556 68474
rect 25504 68410 25556 68416
rect 22744 68400 22796 68406
rect 22744 68342 22796 68348
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21364 3664 21416 3670
rect 20626 3632 20682 3641
rect 21364 3606 21416 3612
rect 20626 3567 20682 3576
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 17052 480 17080 3470
rect 18248 480 18276 3470
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 480 19472 3334
rect 20640 480 20668 3567
rect 21836 480 21864 4966
rect 22756 3602 22784 68342
rect 23020 3800 23072 3806
rect 23020 3742 23072 3748
rect 25318 3768 25374 3777
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 23032 480 23060 3742
rect 25516 3738 25544 68410
rect 25318 3703 25374 3712
rect 25504 3732 25556 3738
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 25332 480 25360 3703
rect 25504 3674 25556 3680
rect 27540 3534 27568 70042
rect 32404 66972 32456 66978
rect 32404 66914 32456 66920
rect 30104 14476 30156 14482
rect 30104 14418 30156 14424
rect 27712 6180 27764 6186
rect 27712 6122 27764 6128
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 26528 480 26556 3470
rect 27724 480 27752 6122
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28920 480 28948 3538
rect 30116 480 30144 14418
rect 32416 6914 32444 66914
rect 32324 6886 32444 6914
rect 31300 3868 31352 3874
rect 31300 3810 31352 3816
rect 31312 480 31340 3810
rect 32324 3670 32352 6886
rect 32312 3664 32364 3670
rect 32312 3606 32364 3612
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 32416 480 32444 3606
rect 34440 3534 34468 70178
rect 37188 68672 37240 68678
rect 37188 68614 37240 68620
rect 35164 68536 35216 68542
rect 35164 68478 35216 68484
rect 34796 6316 34848 6322
rect 34796 6258 34848 6264
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 33612 480 33640 3470
rect 34808 480 34836 6258
rect 35176 3806 35204 68478
rect 35164 3800 35216 3806
rect 35164 3742 35216 3748
rect 35992 3324 36044 3330
rect 35992 3266 36044 3272
rect 36004 480 36032 3266
rect 37200 480 37228 68614
rect 39304 67040 39356 67046
rect 39304 66982 39356 66988
rect 39316 3874 39344 66982
rect 39304 3868 39356 3874
rect 39304 3810 39356 3816
rect 39580 3800 39632 3806
rect 39580 3742 39632 3748
rect 38384 3732 38436 3738
rect 38384 3674 38436 3680
rect 38396 480 38424 3674
rect 39592 480 39620 3742
rect 41340 3398 41368 70246
rect 50344 70168 50396 70174
rect 50344 70110 50396 70116
rect 48228 68740 48280 68746
rect 48228 68682 48280 68688
rect 43444 67108 43496 67114
rect 43444 67050 43496 67056
rect 42800 6384 42852 6390
rect 42800 6326 42852 6332
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 40696 480 40724 3334
<<<<<<< HEAD
rect 42812 2922 42840 6326
rect 43076 3868 43128 3874
rect 43076 3810 43128 3816
rect 41880 2916 41932 2922
rect 41880 2858 41932 2864
rect 42800 2916 42852 2922
rect 42800 2858 42852 2864
rect 41892 480 41920 2858
=======
rect 42812 3194 42840 6326
rect 43076 3868 43128 3874
rect 43076 3810 43128 3816
rect 41880 3188 41932 3194
rect 41880 3130 41932 3136
rect 42800 3188 42852 3194
rect 42800 3130 42852 3136
rect 41892 480 41920 3130
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 43088 480 43116 3810
rect 43456 3738 43484 67050
rect 45376 49020 45428 49026
rect 45376 48962 45428 48968
rect 45388 16574 45416 48962
rect 45388 16546 45508 16574
rect 44272 5092 44324 5098
rect 44272 5034 44324 5040
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 44284 480 44312 5034
rect 45480 480 45508 16546
rect 48240 6914 48268 68682
rect 47872 6886 48268 6914
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 46676 480 46704 3878
rect 47872 480 47900 6886
rect 50356 4962 50384 70110
rect 51724 70032 51776 70038
rect 51724 69974 51776 69980
rect 50988 68332 51040 68338
rect 50988 68274 51040 68280
rect 50344 4956 50396 4962
rect 50344 4898 50396 4904
rect 48964 4208 49016 4214
rect 48964 4150 49016 4156
rect 48976 480 49004 4150
rect 51000 3398 51028 68274
rect 51356 7608 51408 7614
rect 51356 7550 51408 7556
rect 50160 3392 50212 3398
rect 50160 3334 50212 3340
rect 50988 3392 51040 3398
rect 50988 3334 51040 3340
rect 50172 480 50200 3334
rect 51368 480 51396 7550
rect 51736 4214 51764 69974
rect 52552 5160 52604 5166
rect 52552 5102 52604 5108
rect 51724 4208 51776 4214
rect 51724 4150 51776 4156
rect 52564 480 52592 5102
rect 53116 5030 53144 70314
rect 60292 69902 60320 71726
rect 60280 69896 60332 69902
rect 60280 69838 60332 69844
rect 57244 69148 57296 69154
rect 57244 69090 57296 69096
rect 55128 68808 55180 68814
rect 55128 68750 55180 68756
rect 53656 65544 53708 65550
rect 53656 65486 53708 65492
rect 53668 16574 53696 65486
rect 53668 16546 53788 16574
rect 53104 5024 53156 5030
rect 53104 4966 53156 4972
rect 53760 480 53788 16546
rect 55140 6914 55168 68750
rect 54956 6886 55168 6914
rect 54956 480 54984 6886
rect 57256 6254 57284 69090
rect 60660 69086 60688 71726
rect 58624 69080 58676 69086
rect 58624 69022 58676 69028
rect 60648 69080 60700 69086
rect 60648 69022 60700 69028
rect 57244 6248 57296 6254
rect 57244 6190 57296 6196
rect 56048 4956 56100 4962
rect 56048 4898 56100 4904
rect 56060 480 56088 4898
rect 58636 4826 58664 69022
rect 59636 5024 59688 5030
rect 59636 4966 59688 4972
rect 58624 4820 58676 4826
rect 58624 4762 58676 4768
rect 58440 4752 58492 4758
rect 58440 4694 58492 4700
rect 57244 4004 57296 4010
rect 57244 3946 57296 3952
rect 57256 480 57284 3946
rect 58452 480 58480 4694
rect 59648 480 59676 4966
rect 60844 4894 60872 71742
rect 61382 71726 61424 71754
rect 62777 71754 62805 72012
rect 62067 71742 62119 71748
rect 61396 69154 61424 71726
rect 62776 71726 62805 71754
rect 63475 71754 63503 72012
rect 64173 71754 64201 72012
rect 63475 71726 63540 71754
rect 61384 69148 61436 69154
rect 61384 69090 61436 69096
rect 62776 68610 62804 71726
rect 63512 69970 63540 71726
rect 64156 71726 64201 71754
rect 64871 71754 64899 72012
rect 65568 71754 65596 72012
rect 64871 71726 64920 71754
rect 64156 70378 64184 71726
rect 64144 70372 64196 70378
rect 64144 70314 64196 70320
rect 64892 70242 64920 71726
rect 64984 71726 65596 71754
rect 66266 71754 66294 72012
rect 66964 71754 66992 72012
rect 67662 71754 67690 72012
rect 68360 71754 68388 72012
rect 69057 71754 69085 72012
rect 69755 71754 69783 72012
rect 70453 71754 70481 72012
rect 71151 71754 71179 72012
rect 71849 71754 71877 72012
rect 72546 71754 72574 72012
rect 66266 71726 66300 71754
rect 64880 70236 64932 70242
rect 64880 70178 64932 70184
rect 63500 69964 63552 69970
rect 63500 69906 63552 69912
rect 62764 68604 62816 68610
rect 62764 68546 62816 68552
rect 64984 14482 65012 71726
rect 65524 69896 65576 69902
rect 65524 69838 65576 69844
rect 64972 14476 65024 14482
rect 64972 14418 65024 14424
rect 63224 6248 63276 6254
rect 63224 6190 63276 6196
rect 60832 4888 60884 4894
rect 60832 4830 60884 4836
rect 62028 4888 62080 4894
rect 62028 4830 62080 4836
rect 60832 4072 60884 4078
rect 60832 4014 60884 4020
rect 60844 480 60872 4014
rect 62040 480 62068 4830
rect 63236 480 63264 6190
rect 65536 5166 65564 69838
rect 66272 69630 66300 71726
rect 66916 71726 66992 71754
rect 67652 71726 67690 71754
rect 67744 71726 68388 71754
rect 69032 71726 69085 71754
rect 69216 71726 69783 71754
rect 70412 71726 70481 71754
rect 70596 71726 71179 71754
rect 71792 71726 71877 71754
rect 71976 71726 72574 71754
rect 73244 71754 73272 72012
rect 73942 71754 73970 72012
rect 73244 71726 73292 71754
rect 66260 69624 66312 69630
rect 66260 69566 66312 69572
rect 66916 69562 66944 71726
rect 67652 70310 67680 71726
rect 67640 70304 67692 70310
rect 67640 70246 67692 70252
rect 65892 69556 65944 69562
rect 65892 69498 65944 69504
rect 66904 69556 66956 69562
rect 66904 69498 66956 69504
rect 65904 68678 65932 69498
rect 65892 68672 65944 68678
rect 65892 68614 65944 68620
rect 65524 5160 65576 5166
rect 65524 5102 65576 5108
rect 67744 5098 67772 71726
rect 68284 70100 68336 70106
rect 68284 70042 68336 70048
rect 67732 5092 67784 5098
rect 67732 5034 67784 5040
rect 65524 4276 65576 4282
rect 65524 4218 65576 4224
rect 64328 4140 64380 4146
rect 64328 4082 64380 4088
rect 64340 480 64368 4082
rect 65536 480 65564 4218
rect 68296 4214 68324 70042
rect 69032 68746 69060 71726
rect 69020 68740 69072 68746
rect 69020 68682 69072 68688
rect 69216 7614 69244 71726
rect 69664 69080 69716 69086
rect 69664 69022 69716 69028
rect 69204 7608 69256 7614
rect 69204 7550 69256 7556
rect 69112 5568 69164 5574
rect 69112 5510 69164 5516
rect 66720 4208 66772 4214
rect 66720 4150 66772 4156
rect 68284 4208 68336 4214
rect 68284 4150 68336 4156
rect 66732 480 66760 4150
<<<<<<< HEAD
rect 67916 3256 67968 3262
rect 67916 3198 67968 3204
rect 67928 480 67956 3198
=======
rect 67916 3392 67968 3398
rect 67916 3334 67968 3340
rect 67928 480 67956 3334
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 69124 480 69152 5510
rect 69676 4894 69704 69022
rect 70412 68814 70440 71726
rect 70400 68808 70452 68814
rect 70400 68750 70452 68756
rect 70308 7608 70360 7614
rect 70308 7550 70360 7556
rect 69664 4888 69716 4894
rect 69664 4830 69716 4836
rect 70320 480 70348 7550
rect 70596 4758 70624 71726
rect 71792 69086 71820 71726
rect 71780 69080 71832 69086
rect 71780 69022 71832 69028
rect 70584 4752 70636 4758
rect 70584 4694 70636 4700
rect 71976 4282 72004 71726
rect 73264 69154 73292 71726
rect 73908 71726 73970 71754
rect 74640 71754 74668 72012
rect 75338 71754 75366 72012
rect 76035 71754 76063 72012
rect 74640 71726 74672 71754
rect 75338 71726 75408 71754
rect 72424 69148 72476 69154
rect 72424 69090 72476 69096
rect 73252 69148 73304 69154
rect 73252 69090 73304 69096
rect 72436 5574 72464 69090
rect 73908 69086 73936 71726
rect 74644 69154 74672 71726
rect 74632 69148 74684 69154
rect 74632 69090 74684 69096
rect 75380 69086 75408 71726
rect 76024 71726 76063 71754
rect 76733 71754 76761 72012
rect 77431 71754 77459 72012
rect 76733 71726 76788 71754
rect 76024 69154 76052 71726
rect 75736 69148 75788 69154
rect 75736 69090 75788 69096
rect 76012 69148 76064 69154
rect 76012 69090 76064 69096
rect 73068 69080 73120 69086
rect 73068 69022 73120 69028
rect 73896 69080 73948 69086
rect 73896 69022 73948 69028
rect 75368 69080 75420 69086
rect 75368 69022 75420 69028
rect 72424 5568 72476 5574
rect 72424 5510 72476 5516
rect 71964 4276 72016 4282
rect 71964 4218 72016 4224
<<<<<<< HEAD
rect 73080 3398 73108 69022
rect 73804 5160 73856 5166
rect 73804 5102 73856 5108
rect 72608 3392 72660 3398
rect 72608 3334 72660 3340
rect 73068 3392 73120 3398
rect 73068 3334 73120 3340
rect 71504 3188 71556 3194
rect 71504 3130 71556 3136
rect 71516 480 71544 3130
rect 72620 480 72648 3334
=======
rect 71504 3324 71556 3330
rect 71504 3266 71556 3272
rect 71516 480 71544 3266
rect 73080 3262 73108 69022
rect 73804 5160 73856 5166
rect 73804 5102 73856 5108
rect 72608 3256 72660 3262
rect 72608 3198 72660 3204
rect 73068 3256 73120 3262
rect 73068 3198 73120 3204
rect 72620 480 72648 3198
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 73816 480 73844 5102
rect 75748 4214 75776 69090
rect 76760 69086 76788 71726
rect 77404 71726 77459 71754
rect 78129 71754 78157 72012
rect 78827 71754 78855 72012
rect 79524 71754 79552 72012
rect 80222 71754 80250 72012
rect 80920 71754 80948 72012
rect 78129 71726 78168 71754
rect 78827 71726 78904 71754
rect 79524 71726 79916 71754
rect 80222 71726 80284 71754
rect 77116 69148 77168 69154
rect 77116 69090 77168 69096
rect 75828 69080 75880 69086
rect 75828 69022 75880 69028
rect 76748 69080 76800 69086
rect 76748 69022 76800 69028
rect 75840 4282 75868 69022
rect 75828 4276 75880 4282
rect 75828 4218 75880 4224
rect 77128 4214 77156 69090
rect 77404 69086 77432 71726
rect 78140 69222 78168 71726
rect 78128 69216 78180 69222
rect 78128 69158 78180 69164
rect 78876 69154 78904 71726
rect 78864 69148 78916 69154
rect 78864 69090 78916 69096
rect 77208 69080 77260 69086
rect 77208 69022 77260 69028
rect 77392 69080 77444 69086
rect 77392 69022 77444 69028
rect 79324 69080 79376 69086
rect 79324 69022 79376 69028
rect 77220 5098 77248 69022
rect 79336 6526 79364 69022
rect 79324 6520 79376 6526
rect 79324 6462 79376 6468
rect 77392 5296 77444 5302
rect 77392 5238 77444 5244
rect 77208 5092 77260 5098
rect 77208 5034 77260 5040
rect 75736 4208 75788 4214
rect 75736 4150 75788 4156
rect 76196 4208 76248 4214
rect 76196 4150 76248 4156
rect 77116 4208 77168 4214
rect 77116 4150 77168 4156
rect 75000 3256 75052 3262
rect 75000 3198 75052 3204
rect 75012 480 75040 3198
rect 76208 480 76236 4150
rect 77404 480 77432 5238
rect 79888 5234 79916 71726
rect 79968 69148 80020 69154
rect 79968 69090 80020 69096
rect 79980 5438 80008 69090
rect 80256 69086 80284 71726
rect 80900 71726 80948 71754
rect 81618 71754 81646 72012
rect 82316 71754 82344 72012
rect 83013 71754 83041 72012
rect 83711 71754 83739 72012
rect 84409 71754 84437 72012
rect 81618 71726 81664 71754
rect 82316 71726 82400 71754
rect 83013 71726 83044 71754
rect 83711 71726 84056 71754
rect 80900 70174 80928 71726
rect 80888 70168 80940 70174
rect 80888 70110 80940 70116
rect 81636 69630 81664 71726
rect 81624 69624 81676 69630
rect 81624 69566 81676 69572
rect 80244 69080 80296 69086
rect 80244 69022 80296 69028
rect 81348 69080 81400 69086
rect 81348 69022 81400 69028
rect 80888 9104 80940 9110
rect 80888 9046 80940 9052
rect 79968 5432 80020 5438
rect 79968 5374 80020 5380
rect 79876 5228 79928 5234
rect 79876 5170 79928 5176
rect 79692 4276 79744 4282
rect 79692 4218 79744 4224
rect 78588 3188 78640 3194
rect 78588 3130 78640 3136
rect 78600 480 78628 3130
rect 79704 480 79732 4218
rect 80900 480 80928 9046
rect 81360 8974 81388 69022
rect 82372 65686 82400 71726
rect 83016 69086 83044 71726
rect 83464 69216 83516 69222
rect 83464 69158 83516 69164
rect 83004 69080 83056 69086
rect 83004 69022 83056 69028
rect 82360 65680 82412 65686
rect 82360 65622 82412 65628
rect 81348 8968 81400 8974
rect 81348 8910 81400 8916
rect 83476 7682 83504 69158
rect 83464 7676 83516 7682
rect 83464 7618 83516 7624
rect 84028 4826 84056 71726
rect 84396 71726 84437 71754
rect 85107 71754 85135 72012
rect 85805 71754 85833 72012
rect 85107 71726 85160 71754
rect 84396 70242 84424 71726
rect 84384 70236 84436 70242
rect 84384 70178 84436 70184
rect 84108 69080 84160 69086
rect 84108 69022 84160 69028
rect 84120 4894 84148 69022
rect 85132 68406 85160 71726
rect 85776 71726 85833 71754
rect 86502 71754 86530 72012
rect 87200 71890 87228 72012
rect 87156 71862 87228 71890
rect 86502 71726 86540 71754
rect 85776 68474 85804 71726
rect 86224 69624 86276 69630
rect 86224 69566 86276 69572
rect 85764 68468 85816 68474
rect 85764 68410 85816 68416
rect 85120 68400 85172 68406
rect 85120 68342 85172 68348
rect 84476 5364 84528 5370
rect 84476 5306 84528 5312
rect 84108 4888 84160 4894
rect 84108 4830 84160 4836
rect 84016 4820 84068 4826
rect 84016 4762 84068 4768
rect 83280 4208 83332 4214
rect 83280 4150 83332 4156
rect 82084 3120 82136 3126
rect 82084 3062 82136 3068
rect 82096 480 82124 3062
rect 83292 480 83320 4150
rect 84488 480 84516 5306
rect 86236 5098 86264 69566
rect 86512 66978 86540 71726
rect 87156 68542 87184 71862
rect 87898 71754 87926 72012
rect 88596 71890 88624 72012
rect 87340 71726 87926 71754
rect 88536 71862 88624 71890
rect 87144 68536 87196 68542
rect 87144 68478 87196 68484
rect 86500 66972 86552 66978
rect 86500 66914 86552 66920
rect 87340 64874 87368 71726
rect 87604 69080 87656 69086
rect 87604 69022 87656 69028
rect 86972 64846 87368 64874
rect 86972 6186 87000 64846
rect 87616 49026 87644 69022
rect 88536 67046 88564 71862
rect 89294 71754 89322 72012
rect 89991 71890 90019 72012
rect 88628 71726 89322 71754
rect 89824 71862 90019 71890
rect 88524 67040 88576 67046
rect 88524 66982 88576 66988
rect 88628 64874 88656 71726
rect 89824 67114 89852 71862
rect 90689 71754 90717 72012
rect 89916 71726 90717 71754
rect 91387 71754 91415 72012
rect 92085 71754 92113 72012
rect 92783 71890 92811 72012
rect 91387 71726 91416 71754
rect 89812 67108 89864 67114
rect 89812 67050 89864 67056
rect 88352 64846 88656 64874
rect 87604 49020 87656 49026
rect 87604 48962 87656 48968
rect 88352 6322 88380 64846
rect 89916 6390 89944 71726
rect 91388 69086 91416 71726
rect 92032 71726 92113 71754
rect 92492 71862 92811 71890
rect 92032 70038 92060 71726
rect 92020 70032 92072 70038
rect 92020 69974 92072 69980
rect 92492 69902 92520 71862
rect 93480 71754 93508 72012
rect 94178 71754 94206 72012
rect 94876 71754 94904 72012
rect 95574 71754 95602 72012
rect 96272 71754 96300 72012
rect 96969 71754 96997 72012
rect 97667 71754 97695 72012
rect 92584 71726 93508 71754
rect 94148 71726 94206 71754
rect 94332 71726 94904 71754
rect 95528 71726 95602 71754
rect 96264 71726 96300 71754
rect 96724 71726 96997 71754
rect 97644 71726 97695 71754
rect 98000 71800 98052 71806
rect 98365 71754 98393 72012
rect 99063 71806 99091 72012
rect 98000 71742 98052 71748
rect 92480 69896 92532 69902
rect 92480 69838 92532 69844
rect 91376 69080 91428 69086
rect 91376 69022 91428 69028
rect 90364 6520 90416 6526
rect 90364 6462 90416 6468
rect 89904 6384 89956 6390
rect 89904 6326 89956 6332
rect 88340 6316 88392 6322
rect 88340 6258 88392 6264
rect 86960 6180 87012 6186
rect 86960 6122 87012 6128
rect 87972 6180 88024 6186
rect 87972 6122 88024 6128
rect 85764 5092 85816 5098
rect 85764 5034 85816 5040
rect 86224 5092 86276 5098
rect 86224 5034 86276 5040
rect 85776 4214 85804 5034
rect 85764 4208 85816 4214
rect 85764 4150 85816 4156
rect 86868 4208 86920 4214
rect 86868 4150 86920 4156
rect 85672 3052 85724 3058
rect 85672 2994 85724 3000
rect 85684 480 85712 2994
rect 86880 480 86908 4150
rect 87984 480 88012 6122
rect 89168 2984 89220 2990
rect 89168 2926 89220 2932
rect 89180 480 89208 2926
rect 90376 480 90404 6462
rect 92584 4962 92612 71726
rect 94148 69902 94176 71726
rect 93124 69896 93176 69902
rect 93124 69838 93176 69844
rect 94136 69896 94188 69902
rect 94136 69838 94188 69844
rect 93136 5030 93164 69838
rect 94332 64874 94360 71726
rect 95528 70174 95556 71726
rect 95516 70168 95568 70174
rect 95516 70110 95568 70116
rect 94504 69148 94556 69154
rect 94504 69090 94556 69096
rect 93964 64846 94360 64874
rect 93860 7676 93912 7682
rect 93860 7618 93912 7624
rect 93124 5024 93176 5030
rect 93124 4966 93176 4972
rect 92572 4956 92624 4962
rect 92572 4898 92624 4904
rect 91560 4548 91612 4554
rect 91560 4490 91612 4496
rect 91572 480 91600 4490
rect 93872 3482 93900 7618
rect 93964 6254 93992 64846
rect 93952 6248 94004 6254
rect 93952 6190 94004 6196
rect 94516 4554 94544 69090
rect 96264 69086 96292 71726
rect 94596 69080 94648 69086
rect 94596 69022 94648 69028
rect 96252 69080 96304 69086
rect 96252 69022 96304 69028
rect 94608 7614 94636 69022
rect 94596 7608 94648 7614
rect 94596 7550 94648 7556
rect 96724 5166 96752 71726
rect 97644 64874 97672 71726
rect 96816 64846 97672 64874
rect 96816 5302 96844 64846
rect 97448 5432 97500 5438
rect 97448 5374 97500 5380
rect 96804 5296 96856 5302
rect 96804 5238 96856 5244
rect 96712 5160 96764 5166
rect 96712 5102 96764 5108
rect 94504 4548 94556 4554
rect 94504 4490 94556 4496
rect 95148 4208 95200 4214
rect 95148 4150 95200 4156
rect 93872 3454 93992 3482
rect 92756 2916 92808 2922
rect 92756 2858 92808 2864
rect 92768 480 92796 2858
rect 93964 480 93992 3454
rect 95160 480 95188 4150
rect 96252 2848 96304 2854
rect 96252 2790 96304 2796
rect 96264 480 96292 2790
rect 97460 480 97488 5374
rect 98012 5370 98040 71742
rect 98104 71726 98393 71754
rect 99051 71800 99103 71806
rect 99761 71754 99789 72012
rect 100458 71754 100486 72012
rect 99051 71742 99103 71748
rect 99760 71726 99789 71754
rect 100404 71726 100486 71754
rect 100760 71800 100812 71806
rect 101156 71754 101184 72012
rect 101854 71806 101882 72012
rect 100760 71742 100812 71748
rect 98104 9110 98132 71726
rect 99760 69086 99788 71726
rect 100404 69154 100432 71726
rect 100668 69624 100720 69630
rect 100668 69566 100720 69572
rect 100392 69148 100444 69154
rect 100392 69090 100444 69096
rect 98644 69080 98696 69086
rect 98644 69022 98696 69028
rect 99748 69080 99800 69086
rect 99748 69022 99800 69028
rect 98092 9104 98144 9110
rect 98092 9046 98144 9052
rect 98656 6186 98684 69022
rect 100680 6914 100708 69566
rect 100312 6886 100708 6914
rect 98644 6180 98696 6186
rect 98644 6122 98696 6128
rect 98644 5568 98696 5574
rect 98644 5510 98696 5516
rect 98000 5364 98052 5370
rect 98000 5306 98052 5312
rect 98656 480 98684 5510
<<<<<<< HEAD
rect 100312 2854 100340 6886
=======
rect 99852 598 100064 626
rect 99852 480 99880 598
rect 100036 490 100064 598
rect 100312 490 100340 6886
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 100772 5574 100800 71742
rect 100956 71726 101184 71754
rect 101842 71800 101894 71806
rect 102552 71754 102580 72012
rect 101842 71742 101894 71748
rect 102152 71726 102580 71754
rect 103250 71754 103278 72012
rect 103947 71754 103975 72012
rect 104645 71754 104673 72012
rect 105343 71754 105371 72012
rect 106041 71754 106069 72012
rect 106739 71754 106767 72012
rect 107436 71754 107464 72012
rect 108134 71890 108162 72012
rect 103250 71726 103284 71754
rect 103947 71726 104020 71754
rect 104645 71726 104756 71754
rect 105343 71726 105400 71754
rect 106041 71726 106228 71754
rect 106739 71726 106780 71754
rect 100760 5568 100812 5574
rect 100760 5510 100812 5516
rect 100956 4214 100984 71726
rect 102152 16574 102180 71726
rect 103256 69902 103284 71726
rect 103428 70100 103480 70106
rect 103428 70042 103480 70048
rect 103244 69896 103296 69902
rect 103244 69838 103296 69844
rect 102152 16546 102272 16574
rect 101036 5228 101088 5234
rect 101036 5170 101088 5176
rect 100944 4208 100996 4214
rect 100944 4150 100996 4156
<<<<<<< HEAD
rect 99840 2848 99892 2854
rect 99840 2790 99892 2796
rect 100300 2848 100352 2854
rect 100300 2790 100352 2796
rect 99852 480 99880 2790
rect 101048 480 101076 5170
rect 102244 480 102272 16546
rect 103440 6914 103468 70042
rect 103992 69086 104020 71726
rect 104164 69896 104216 69902
rect 104164 69838 104216 69844
rect 103980 69080 104032 69086
rect 103980 69022 104032 69028
rect 104176 14142 104204 69838
rect 104164 14136 104216 14142
rect 104164 14078 104216 14084
rect 104532 8968 104584 8974
rect 104532 8910 104584 8916
rect 103348 6886 103468 6914
rect 103348 480 103376 6886
rect 104544 480 104572 8910
rect 104728 5574 104756 71726
rect 105372 69086 105400 71726
rect 104808 69080 104860 69086
rect 104808 69022 104860 69028
rect 105360 69080 105412 69086
rect 105360 69022 105412 69028
rect 106096 69080 106148 69086
rect 106096 69022 106148 69028
rect 104716 5568 104768 5574
rect 104716 5510 104768 5516
rect 104820 4214 104848 69022
rect 105728 14136 105780 14142
rect 105728 14078 105780 14084
rect 104808 4208 104860 4214
rect 104808 4150 104860 4156
rect 105740 480 105768 14078
rect 106108 7614 106136 69022
rect 106096 7608 106148 7614
rect 106096 7550 106148 7556
rect 106200 4962 106228 71726
rect 106752 70174 106780 71726
rect 107396 71726 107464 71754
rect 107672 71862 108162 71890
rect 106740 70168 106792 70174
rect 106740 70110 106792 70116
rect 107396 66910 107424 71726
rect 107476 70100 107528 70106
rect 107476 70042 107528 70048
rect 107384 66904 107436 66910
rect 107384 66846 107436 66852
rect 107488 64874 107516 70042
rect 107568 69964 107620 69970
rect 107568 69906 107620 69912
rect 107580 69714 107608 69906
rect 107672 69834 107700 71862
rect 108832 71754 108860 72012
rect 107764 71726 108860 71754
rect 109132 71800 109184 71806
rect 109530 71754 109558 72012
rect 110228 71806 110256 72012
rect 109132 71742 109184 71748
rect 107660 69828 107712 69834
rect 107660 69770 107712 69776
rect 107580 69686 107700 69714
rect 107488 64846 107608 64874
rect 106188 4956 106240 4962
rect 106188 4898 106240 4904
rect 107580 3534 107608 64846
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 107672 3482 107700 69686
rect 107764 4010 107792 71726
rect 107752 4004 107804 4010
rect 107752 3946 107804 3952
rect 109144 3602 109172 71742
rect 109236 71726 109558 71754
rect 110216 71800 110268 71806
rect 110925 71754 110953 72012
rect 111623 71754 111651 72012
rect 112321 71754 112349 72012
rect 113019 71754 113047 72012
rect 113717 71754 113745 72012
rect 114414 71754 114442 72012
rect 110216 71742 110268 71748
rect 110524 71726 110953 71754
rect 110984 71726 111651 71754
rect 111904 71726 112349 71754
rect 112456 71726 113047 71754
rect 113284 71726 113745 71754
rect 114388 71726 114442 71754
rect 114560 71800 114612 71806
rect 114560 71742 114612 71748
rect 115112 71754 115140 72012
rect 115810 71806 115838 72012
rect 115798 71800 115850 71806
rect 109236 4282 109264 71726
rect 109224 4276 109276 4282
rect 109224 4218 109276 4224
rect 109316 4208 109368 4214
rect 109316 4150 109368 4156
rect 109132 3596 109184 3602
rect 109132 3538 109184 3544
rect 106936 480 106964 3470
rect 107672 3454 108160 3482
rect 108132 480 108160 3454
rect 109328 480 109356 4150
rect 110524 3670 110552 71726
rect 110984 64874 111012 71726
rect 111708 69828 111760 69834
rect 111708 69770 111760 69776
rect 110616 64846 111012 64874
rect 110616 3738 110644 64846
rect 111616 5092 111668 5098
rect 111616 5034 111668 5040
rect 110604 3732 110656 3738
rect 110604 3674 110656 3680
rect 110512 3664 110564 3670
rect 110512 3606 110564 3612
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 110524 480 110552 3470
rect 111628 480 111656 5034
rect 111720 3534 111748 69770
rect 111800 69284 111852 69290
rect 111800 69226 111852 69232
rect 111812 68338 111840 69226
rect 111800 68332 111852 68338
rect 111800 68274 111852 68280
rect 111904 3806 111932 71726
rect 112456 64874 112484 71726
rect 111996 64846 112484 64874
rect 111996 3874 112024 64846
rect 112812 5568 112864 5574
rect 112812 5510 112864 5516
rect 111984 3868 112036 3874
rect 111984 3810 112036 3816
rect 111892 3800 111944 3806
rect 111892 3742 111944 3748
rect 111708 3528 111760 3534
rect 111708 3470 111760 3476
rect 112824 480 112852 5510
rect 113284 3534 113312 71726
rect 114388 69290 114416 71726
rect 114468 69964 114520 69970
rect 114468 69906 114520 69912
rect 114376 69284 114428 69290
rect 114376 69226 114428 69232
rect 113272 3528 113324 3534
rect 113272 3470 113324 3476
rect 114480 3330 114508 69906
rect 114572 3466 114600 71742
rect 115112 71726 115152 71754
rect 115798 71742 115850 71748
rect 116032 71800 116084 71806
rect 116508 71754 116536 72012
rect 117206 71806 117234 72012
rect 116032 71742 116084 71748
rect 114652 65680 114704 65686
rect 114652 65622 114704 65628
rect 114664 16574 114692 65622
rect 115124 65550 115152 71726
rect 115112 65544 115164 65550
rect 115112 65486 115164 65492
rect 114664 16546 115244 16574
rect 114560 3460 114612 3466
rect 114560 3402 114612 3408
rect 114008 3324 114060 3330
rect 114008 3266 114060 3272
rect 114468 3324 114520 3330
rect 114468 3266 114520 3272
rect 114020 480 114048 3266
rect 115216 480 115244 16546
rect 116044 4146 116072 71742
rect 116136 71726 116536 71754
rect 117194 71800 117246 71806
rect 117194 71742 117246 71748
rect 117320 71800 117372 71806
rect 117903 71754 117931 72012
rect 118601 71806 118629 72012
rect 117320 71742 117372 71748
rect 116032 4140 116084 4146
rect 116032 4082 116084 4088
rect 116136 4078 116164 71726
rect 116400 7608 116452 7614
rect 116400 7550 116452 7556
rect 116124 4072 116176 4078
rect 116124 4014 116176 4020
rect 116412 480 116440 7550
rect 116492 4956 116544 4962
rect 116492 4898 116544 4904
rect 116504 2922 116532 4898
rect 117332 3262 117360 71742
rect 117424 71726 117931 71754
rect 118589 71800 118641 71806
rect 118589 71742 118641 71748
rect 118792 71800 118844 71806
rect 119299 71754 119327 72012
rect 119997 71806 120025 72012
rect 118792 71742 118844 71748
rect 117424 3398 117452 71726
rect 118804 6914 118832 71742
rect 118712 6886 118832 6914
rect 118988 71726 119327 71754
rect 119985 71800 120037 71806
rect 119985 71742 120037 71748
rect 120172 71800 120224 71806
rect 120695 71754 120723 72012
rect 121392 71806 121420 72012
rect 120172 71742 120224 71748
rect 117412 3392 117464 3398
rect 117412 3334 117464 3340
rect 117320 3256 117372 3262
rect 117320 3198 117372 3204
rect 118712 3194 118740 6886
rect 118792 4888 118844 4894
rect 118792 4830 118844 4836
rect 118700 3188 118752 3194
rect 118700 3130 118752 3136
rect 117596 3052 117648 3058
rect 117596 2994 117648 3000
rect 116492 2916 116544 2922
rect 116492 2858 116544 2864
rect 117608 480 117636 2994
rect 118804 480 118832 4830
rect 118988 3534 119016 71726
rect 119344 70236 119396 70242
rect 119344 70178 119396 70184
rect 118976 3528 119028 3534
rect 118976 3470 119028 3476
rect 119356 3058 119384 70178
rect 119344 3052 119396 3058
rect 119344 2994 119396 3000
rect 120184 2990 120212 71742
rect 120276 71726 120723 71754
rect 121380 71800 121432 71806
rect 122090 71754 122118 72012
rect 122788 71754 122816 72012
rect 123486 71754 123514 72012
rect 124184 71754 124212 72012
rect 124881 71754 124909 72012
rect 121380 71742 121432 71748
rect 121564 71726 122118 71754
rect 122208 71726 122816 71754
rect 122944 71726 123514 71754
rect 124140 71726 124212 71754
rect 124876 71726 124909 71754
rect 125579 71754 125607 72012
rect 126277 71754 126305 72012
rect 125579 71726 125640 71754
rect 120276 3126 120304 71726
rect 121368 70304 121420 70310
rect 121368 70246 121420 70252
rect 121380 6914 121408 70246
rect 121104 6886 121408 6914
rect 120264 3120 120316 3126
rect 120264 3062 120316 3068
rect 120172 2984 120224 2990
rect 120172 2926 120224 2932
rect 119896 2916 119948 2922
rect 119896 2858 119948 2864
rect 119908 480 119936 2858
rect 121104 480 121132 6886
rect 121564 3330 121592 71726
rect 122208 64874 122236 71726
rect 122840 70168 122892 70174
rect 122840 70110 122892 70116
rect 121656 64846 122236 64874
rect 121656 3466 121684 64846
rect 122288 4820 122340 4826
rect 122288 4762 122340 4768
rect 121644 3460 121696 3466
rect 121644 3402 121696 3408
rect 121552 3324 121604 3330
rect 121552 3266 121604 3272
rect 122300 480 122328 4762
rect 122852 2666 122880 70110
rect 122944 2854 122972 71726
rect 124140 69902 124168 71726
rect 124876 70038 124904 71726
rect 125612 70106 125640 71726
rect 126256 71726 126305 71754
rect 126975 71754 127003 72012
rect 127673 71754 127701 72012
rect 126975 71726 127020 71754
rect 125600 70100 125652 70106
rect 125600 70042 125652 70048
rect 124864 70032 124916 70038
rect 124864 69974 124916 69980
rect 124128 69896 124180 69902
rect 124128 69838 124180 69844
rect 126256 69834 126284 71726
rect 126992 69970 127020 71726
rect 127636 71726 127701 71754
rect 128370 71754 128398 72012
rect 129068 71754 129096 72012
rect 128370 71726 128400 71754
rect 127636 70242 127664 71726
rect 128372 70310 128400 71726
rect 129016 71726 129096 71754
rect 129766 71754 129794 72012
rect 130464 71754 130492 72012
rect 131162 71754 131190 72012
rect 131859 71754 131887 72012
rect 129766 71726 129872 71754
rect 130464 71726 130516 71754
rect 128360 70304 128412 70310
rect 128360 70246 128412 70252
rect 127624 70236 127676 70242
rect 127624 70178 127676 70184
rect 126980 69964 127032 69970
rect 126980 69906 127032 69912
rect 126244 69828 126296 69834
rect 126244 69770 126296 69776
rect 126888 69420 126940 69426
rect 126888 69362 126940 69368
rect 125508 69080 125560 69086
rect 125508 69022 125560 69028
rect 125520 3534 125548 69022
rect 126900 3534 126928 69362
rect 129016 69086 129044 71726
rect 129648 69828 129700 69834
rect 129648 69770 129700 69776
rect 129004 69080 129056 69086
rect 129004 69022 129056 69028
rect 129660 16574 129688 69770
rect 129384 16546 129688 16574
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 122932 2848 122984 2854
rect 122932 2790 122984 2796
rect 122852 2638 123524 2666
rect 123496 480 123524 2638
rect 124692 480 124720 3470
rect 125888 480 125916 3470
rect 128176 3460 128228 3466
rect 128176 3402 128228 3408
rect 126980 3120 127032 3126
rect 126980 3062 127032 3068
rect 126992 480 127020 3062
rect 128188 480 128216 3402
rect 129384 480 129412 16546
rect 129648 9240 129700 9246
rect 129648 9182 129700 9188
rect 129660 3126 129688 9182
rect 129844 3505 129872 71726
rect 130488 69766 130516 71726
rect 131132 71726 131190 71754
rect 131224 71726 131887 71754
rect 132557 71754 132585 72012
rect 133255 71754 133283 72012
rect 133953 71754 133981 72012
rect 134651 71754 134679 72012
rect 132557 71726 132632 71754
rect 131028 69896 131080 69902
rect 131028 69838 131080 69844
rect 130476 69760 130528 69766
rect 130476 69702 130528 69708
rect 131040 3534 131068 69838
rect 131132 3641 131160 71726
rect 131224 3777 131252 71726
rect 131764 3868 131816 3874
rect 131764 3810 131816 3816
rect 131210 3768 131266 3777
rect 131210 3703 131266 3712
rect 131118 3632 131174 3641
rect 131118 3567 131174 3576
rect 130568 3528 130620 3534
rect 129830 3496 129886 3505
rect 130568 3470 130620 3476
rect 131028 3528 131080 3534
rect 131028 3470 131080 3476
rect 129830 3431 129886 3440
rect 129648 3120 129700 3126
rect 129648 3062 129700 3068
rect 130580 480 130608 3470
rect 131776 480 131804 3810
rect 132604 3369 132632 71726
rect 133248 71726 133283 71754
rect 133892 71726 133981 71754
rect 134628 71726 134679 71754
rect 135348 71754 135376 72012
rect 136046 71754 136074 72012
rect 135348 71726 135392 71754
rect 133248 69698 133276 71726
rect 133236 69692 133288 69698
rect 133236 69634 133288 69640
rect 133892 69426 133920 71726
rect 134628 69834 134656 71726
rect 135168 70032 135220 70038
rect 135168 69974 135220 69980
rect 134616 69828 134668 69834
rect 134616 69770 134668 69776
rect 133880 69420 133932 69426
rect 133880 69362 133932 69368
rect 133788 69080 133840 69086
rect 133788 69022 133840 69028
rect 133800 3534 133828 69022
rect 134524 68332 134576 68338
rect 134524 68274 134576 68280
rect 134536 3534 134564 68274
rect 132960 3528 133012 3534
rect 132960 3470 133012 3476
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 134524 3528 134576 3534
rect 134524 3470 134576 3476
rect 132590 3360 132646 3369
rect 132590 3295 132646 3304
rect 132972 480 133000 3470
rect 135180 3466 135208 69974
rect 135364 69086 135392 71726
rect 135456 71726 136074 71754
rect 135352 69080 135404 69086
rect 135352 69022 135404 69028
rect 135260 3800 135312 3806
rect 135260 3742 135312 3748
rect 134156 3460 134208 3466
rect 134156 3402 134208 3408
rect 135168 3460 135220 3466
rect 135168 3402 135220 3408
rect 134168 480 134196 3402
rect 135272 480 135300 3742
rect 135456 2922 135484 71726
rect 136744 69086 136772 72012
rect 137442 71754 137470 72012
rect 138140 71754 138168 72012
rect 137442 71726 137784 71754
rect 136732 69080 136784 69086
rect 136732 69022 136784 69028
rect 137756 4146 137784 71726
rect 138124 71726 138168 71754
rect 138837 71754 138865 72012
rect 139535 71754 139563 72012
rect 140233 71754 140261 72012
rect 140931 71754 140959 72012
rect 141629 71754 141657 72012
rect 142326 71754 142354 72012
rect 143024 71754 143052 72012
rect 143722 71754 143750 72012
rect 144420 71754 144448 72012
rect 145118 71754 145146 72012
rect 138837 71726 139256 71754
rect 139535 71726 139624 71754
rect 140233 71726 140636 71754
rect 140931 71726 141004 71754
rect 141629 71726 141924 71754
rect 142326 71726 142384 71754
rect 143024 71726 143396 71754
rect 143722 71726 143764 71754
rect 144420 71726 144776 71754
rect 137928 70168 137980 70174
rect 137928 70110 137980 70116
rect 137836 69080 137888 69086
rect 137836 69022 137888 69028
rect 137744 4140 137796 4146
rect 137744 4082 137796 4088
rect 137848 3602 137876 69022
rect 137836 3596 137888 3602
rect 137836 3538 137888 3544
rect 137940 3482 137968 70110
rect 138124 69086 138152 71726
rect 138112 69080 138164 69086
rect 138112 69022 138164 69028
rect 139228 3670 139256 71726
rect 139596 69086 139624 71726
rect 139308 69080 139360 69086
rect 139308 69022 139360 69028
rect 139584 69080 139636 69086
rect 139584 69022 139636 69028
rect 139216 3664 139268 3670
rect 139216 3606 139268 3612
rect 139320 3534 139348 69022
rect 140608 3942 140636 71726
rect 140976 69086 141004 71726
rect 140688 69080 140740 69086
rect 140688 69022 140740 69028
rect 140964 69080 141016 69086
rect 140964 69022 141016 69028
rect 140596 3936 140648 3942
rect 140596 3878 140648 3884
rect 140700 3670 140728 69022
rect 141896 6186 141924 71726
rect 141976 70304 142028 70310
rect 141976 70246 142028 70252
rect 141884 6180 141936 6186
rect 141884 6122 141936 6128
rect 140688 3664 140740 3670
rect 140688 3606 140740 3612
rect 140044 3596 140096 3602
rect 140044 3538 140096 3544
rect 137664 3454 137968 3482
rect 139308 3528 139360 3534
rect 139308 3470 139360 3476
rect 135444 2916 135496 2922
rect 135444 2858 135496 2864
rect 136456 2916 136508 2922
rect 136456 2858 136508 2864
rect 136468 480 136496 2858
rect 137664 480 137692 3454
rect 138846 3360 138902 3369
rect 138846 3295 138902 3304
rect 138860 480 138888 3295
rect 140056 480 140084 3538
rect 141988 3058 142016 70246
rect 142356 69086 142384 71726
rect 142068 69080 142120 69086
rect 142068 69022 142120 69028
rect 142344 69080 142396 69086
rect 142344 69022 142396 69028
rect 142080 3738 142108 69022
rect 143368 4554 143396 71726
rect 143736 69086 143764 71726
rect 143448 69080 143500 69086
rect 143448 69022 143500 69028
rect 143724 69080 143776 69086
rect 143724 69022 143776 69028
rect 144644 69080 144696 69086
rect 144644 69022 144696 69028
rect 143356 4548 143408 4554
rect 143356 4490 143408 4496
rect 143460 4486 143488 69022
rect 144656 16574 144684 69022
rect 144564 16546 144684 16574
rect 144564 4622 144592 16546
rect 144748 11778 144776 71726
rect 145116 71726 145146 71754
rect 145815 71754 145843 72012
rect 146513 71754 146541 72012
rect 145815 71726 146248 71754
rect 144828 70236 144880 70242
rect 144828 70178 144880 70184
rect 144656 11750 144776 11778
rect 144656 4690 144684 11750
rect 144840 6914 144868 70178
rect 145116 69086 145144 71726
rect 145104 69080 145156 69086
rect 145104 69022 145156 69028
rect 146116 69080 146168 69086
rect 146116 69022 146168 69028
rect 144748 6886 144868 6914
rect 144644 4684 144696 4690
rect 144644 4626 144696 4632
rect 144552 4616 144604 4622
rect 144552 4558 144604 4564
rect 143448 4480 143500 4486
rect 143448 4422 143500 4428
rect 143540 4140 143592 4146
rect 143540 4082 143592 4088
rect 142068 3732 142120 3738
rect 142068 3674 142120 3680
rect 142434 3496 142490 3505
rect 142434 3431 142490 3440
rect 141240 3052 141292 3058
rect 141240 2994 141292 3000
rect 141976 3052 142028 3058
rect 141976 2994 142028 3000
rect 141252 480 141280 2994
rect 142448 480 142476 3431
rect 143552 480 143580 4082
rect 144748 480 144776 6886
rect 146128 4758 146156 69022
rect 146220 5506 146248 71726
rect 146496 71726 146541 71754
rect 147211 71754 147239 72012
rect 147909 71754 147937 72012
rect 148607 71754 148635 72012
rect 149304 71754 149332 72012
rect 150002 71754 150030 72012
rect 150700 71754 150728 72012
rect 151398 71754 151426 72012
rect 152096 71754 152124 72012
rect 152793 71754 152821 72012
rect 153491 71754 153519 72012
rect 147211 71726 147536 71754
rect 147909 71726 147996 71754
rect 148607 71726 148824 71754
rect 149304 71726 149376 71754
rect 150002 71726 150388 71754
rect 150700 71726 150756 71754
rect 151398 71726 151676 71754
rect 152096 71726 152136 71754
rect 152793 71726 153148 71754
rect 146496 69086 146524 71726
rect 146484 69080 146536 69086
rect 146484 69022 146536 69028
rect 146208 5500 146260 5506
rect 146208 5442 146260 5448
rect 147508 5370 147536 71726
rect 147968 69086 147996 71726
rect 147588 69080 147640 69086
rect 147588 69022 147640 69028
rect 147956 69080 148008 69086
rect 147956 69022 148008 69028
rect 147600 5438 147628 69022
rect 147588 5432 147640 5438
rect 147588 5374 147640 5380
rect 147496 5364 147548 5370
rect 147496 5306 147548 5312
rect 148796 5234 148824 71726
rect 148968 70372 149020 70378
rect 148968 70314 149020 70320
rect 148876 69080 148928 69086
rect 148876 69022 148928 69028
rect 148888 5302 148916 69022
rect 148876 5296 148928 5302
rect 148876 5238 148928 5244
rect 148784 5228 148836 5234
rect 148784 5170 148836 5176
rect 146116 4752 146168 4758
rect 146116 4694 146168 4700
rect 148980 3534 149008 70314
rect 149348 69086 149376 71726
rect 149336 69080 149388 69086
rect 149336 69022 149388 69028
rect 150256 69080 150308 69086
rect 150256 69022 150308 69028
rect 150268 5166 150296 69022
rect 150256 5160 150308 5166
rect 150256 5102 150308 5108
rect 150360 5098 150388 71726
rect 150728 69086 150756 71726
rect 150716 69080 150768 69086
rect 150716 69022 150768 69028
rect 150348 5092 150400 5098
rect 150348 5034 150400 5040
rect 151648 4962 151676 71726
rect 152108 69086 152136 71726
rect 151728 69080 151780 69086
rect 151728 69022 151780 69028
rect 152096 69080 152148 69086
rect 152096 69022 152148 69028
rect 153016 69080 153068 69086
rect 153016 69022 153068 69028
rect 151740 5030 151768 69022
rect 151728 5024 151780 5030
rect 151728 4966 151780 4972
rect 151636 4956 151688 4962
rect 151636 4898 151688 4904
rect 153028 4894 153056 69022
rect 153016 4888 153068 4894
rect 153016 4830 153068 4836
rect 153120 4826 153148 71726
rect 153488 71726 153519 71754
rect 154189 71754 154217 72012
rect 154887 71754 154915 72012
rect 154189 71726 154252 71754
rect 153488 69086 153516 71726
rect 154224 69834 154252 71726
rect 154868 71726 154915 71754
rect 155585 71754 155613 72012
rect 156282 71754 156310 72012
rect 156980 71754 157008 72012
rect 157678 71754 157706 72012
rect 158376 71754 158404 72012
rect 159074 71754 159102 72012
rect 159771 71754 159799 72012
rect 160469 71754 160497 72012
rect 161167 71754 161195 72012
rect 161865 71754 161893 72012
rect 155585 71726 155816 71754
rect 156282 71726 156368 71754
rect 156980 71726 157288 71754
rect 157678 71726 157748 71754
rect 158376 71726 158668 71754
rect 159074 71726 159128 71754
rect 159771 71726 160048 71754
rect 160469 71726 160508 71754
rect 161167 71726 161336 71754
rect 154212 69828 154264 69834
rect 154212 69770 154264 69776
rect 154868 69426 154896 71726
rect 154856 69420 154908 69426
rect 154856 69362 154908 69368
rect 153476 69080 153528 69086
rect 153476 69022 153528 69028
rect 154488 69080 154540 69086
rect 154488 69022 154540 69028
rect 153108 4820 153160 4826
rect 153108 4762 153160 4768
rect 154500 4282 154528 69022
rect 155788 6662 155816 71726
rect 155868 69624 155920 69630
rect 155868 69566 155920 69572
rect 155776 6656 155828 6662
rect 155776 6598 155828 6604
rect 154488 4276 154540 4282
rect 154488 4218 154540 4224
rect 154212 3664 154264 3670
rect 154212 3606 154264 3612
rect 150624 3596 150676 3602
rect 150624 3538 150676 3544
rect 153016 3596 153068 3602
rect 153016 3538 153068 3544
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 145932 3460 145984 3466
rect 145932 3402 145984 3408
rect 145944 480 145972 3402
rect 147140 480 147168 3470
rect 148336 480 148364 3470
rect 149532 480 149560 3470
rect 150636 480 150664 3538
rect 151820 3324 151872 3330
rect 151820 3266 151872 3272
rect 151832 480 151860 3266
rect 153028 480 153056 3538
rect 154224 480 154252 3606
rect 155880 3194 155908 69566
rect 156340 69358 156368 71726
rect 156328 69352 156380 69358
rect 156328 69294 156380 69300
rect 157260 6594 157288 71726
rect 157720 69562 157748 71726
rect 157708 69556 157760 69562
rect 157708 69498 157760 69504
rect 158640 10606 158668 71726
rect 159100 69086 159128 71726
rect 159088 69080 159140 69086
rect 159088 69022 159140 69028
rect 159916 69080 159968 69086
rect 159916 69022 159968 69028
rect 158628 10600 158680 10606
rect 158628 10542 158680 10548
rect 159928 10538 159956 69022
rect 159916 10532 159968 10538
rect 159916 10474 159968 10480
rect 157248 6588 157300 6594
rect 157248 6530 157300 6536
rect 160020 6526 160048 71726
rect 160480 69086 160508 71726
rect 160468 69080 160520 69086
rect 160468 69022 160520 69028
rect 160744 12096 160796 12102
rect 160744 12038 160796 12044
rect 160008 6520 160060 6526
rect 160008 6462 160060 6468
rect 157800 3936 157852 3942
rect 157800 3878 157852 3884
rect 158904 3936 158956 3942
rect 158904 3878 158956 3884
rect 156604 3664 156656 3670
rect 156604 3606 156656 3612
rect 155408 3188 155460 3194
rect 155408 3130 155460 3136
rect 155868 3188 155920 3194
rect 155868 3130 155920 3136
rect 155420 480 155448 3130
rect 156616 480 156644 3606
rect 157812 480 157840 3878
rect 158916 480 158944 3878
rect 160100 3732 160152 3738
rect 160100 3674 160152 3680
rect 160112 480 160140 3674
rect 160756 3330 160784 12038
rect 161308 10402 161336 71726
rect 161860 71726 161893 71754
rect 162563 71754 162591 72012
rect 163260 71754 163288 72012
rect 162563 71726 162808 71754
rect 161860 69086 161888 71726
rect 161388 69080 161440 69086
rect 161388 69022 161440 69028
rect 161848 69080 161900 69086
rect 161848 69022 161900 69028
rect 162676 69080 162728 69086
rect 162676 69022 162728 69028
rect 161400 10470 161428 69022
rect 162124 18624 162176 18630
rect 162124 18566 162176 18572
rect 161388 10464 161440 10470
rect 161388 10406 161440 10412
rect 161296 10396 161348 10402
rect 161296 10338 161348 10344
rect 162136 3874 162164 18566
rect 162688 12034 162716 69022
rect 162676 12028 162728 12034
rect 162676 11970 162728 11976
rect 162492 10668 162544 10674
rect 162492 10610 162544 10616
rect 162124 3868 162176 3874
rect 162124 3810 162176 3816
rect 161296 3392 161348 3398
rect 161296 3334 161348 3340
rect 160744 3324 160796 3330
rect 160744 3266 160796 3272
rect 161308 480 161336 3334
rect 162504 480 162532 10610
rect 162780 10334 162808 71726
rect 163240 71726 163288 71754
rect 163958 71754 163986 72012
rect 164656 71754 164684 72012
rect 165354 71754 165382 72012
rect 166052 71754 166080 72012
rect 166749 71754 166777 72012
rect 167447 71754 167475 72012
rect 168145 71754 168173 72012
rect 168843 71754 168871 72012
rect 169541 71754 169569 72012
rect 170238 71754 170266 72012
rect 163958 71726 164004 71754
rect 164656 71726 164740 71754
rect 165354 71726 165568 71754
rect 166052 71726 166120 71754
rect 166749 71726 166948 71754
rect 167447 71726 167500 71754
rect 168145 71726 168236 71754
rect 168843 71726 168880 71754
rect 169541 71726 169616 71754
rect 163240 69290 163268 71726
rect 163976 70106 164004 71726
rect 163964 70100 164016 70106
rect 163964 70042 164016 70048
rect 164712 69494 164740 71726
rect 164700 69488 164752 69494
rect 164700 69430 164752 69436
rect 163228 69284 163280 69290
rect 163228 69226 163280 69232
rect 164148 15972 164200 15978
rect 164148 15914 164200 15920
rect 162768 10328 162820 10334
rect 162768 10270 162820 10276
rect 164160 3398 164188 15914
rect 165540 11898 165568 71726
rect 166092 69086 166120 71726
rect 166080 69080 166132 69086
rect 166080 69022 166132 69028
rect 166816 69080 166868 69086
rect 166816 69022 166868 69028
rect 165528 11892 165580 11898
rect 165528 11834 165580 11840
rect 166828 6390 166856 69022
rect 166816 6384 166868 6390
rect 166816 6326 166868 6332
rect 166920 6322 166948 71726
rect 167472 69086 167500 71726
rect 167460 69080 167512 69086
rect 167460 69022 167512 69028
rect 167184 6452 167236 6458
rect 167184 6394 167236 6400
rect 166908 6316 166960 6322
rect 166908 6258 166960 6264
rect 164884 6180 164936 6186
rect 164884 6122 164936 6128
rect 163688 3392 163740 3398
rect 163688 3334 163740 3340
rect 164148 3392 164200 3398
rect 164148 3334 164200 3340
rect 163700 480 163728 3334
rect 164896 480 164924 6122
rect 166080 3188 166132 3194
rect 166080 3130 166132 3136
rect 166092 480 166120 3130
rect 167196 480 167224 6394
rect 168208 6186 168236 71726
rect 168852 69086 168880 71726
rect 168288 69080 168340 69086
rect 168288 69022 168340 69028
rect 168840 69080 168892 69086
rect 168840 69022 168892 69028
rect 168300 6254 168328 69022
rect 169588 13530 169616 71726
rect 170232 71726 170266 71754
rect 170936 71754 170964 72012
rect 171634 71754 171662 72012
rect 170936 71726 171088 71754
rect 170232 69086 170260 71726
rect 169668 69080 169720 69086
rect 169668 69022 169720 69028
rect 170220 69080 170272 69086
rect 170220 69022 170272 69028
rect 170956 69080 171008 69086
rect 170956 69022 171008 69028
rect 169576 13524 169628 13530
rect 169576 13466 169628 13472
rect 169680 12306 169708 69022
rect 170968 14754 170996 69022
rect 170956 14748 171008 14754
rect 170956 14690 171008 14696
rect 170404 14544 170456 14550
rect 170404 14486 170456 14492
rect 169668 12300 169720 12306
rect 169668 12242 169720 12248
rect 169576 12164 169628 12170
rect 169576 12106 169628 12112
rect 168288 6248 168340 6254
rect 168288 6190 168340 6196
rect 168196 6180 168248 6186
rect 168196 6122 168248 6128
rect 168380 4480 168432 4486
rect 168380 4422 168432 4428
rect 168392 480 168420 4422
rect 169588 480 169616 12106
rect 170416 3194 170444 14486
rect 171060 12238 171088 71726
rect 171612 71726 171662 71754
rect 172332 71754 172360 72012
rect 173030 71754 173058 72012
rect 173727 71754 173755 72012
rect 174425 71754 174453 72012
rect 175123 71754 175151 72012
rect 175821 71754 175849 72012
rect 176519 71754 176547 72012
rect 177216 71754 177244 72012
rect 177914 71754 177942 72012
rect 178612 71754 178640 72012
rect 172332 71726 172376 71754
rect 173030 71726 173112 71754
rect 173727 71726 173756 71754
rect 174425 71726 174492 71754
rect 175123 71726 175228 71754
rect 175821 71726 175872 71754
rect 176519 71726 176608 71754
rect 177216 71726 177252 71754
rect 171612 69086 171640 71726
rect 171600 69080 171652 69086
rect 171600 69022 171652 69028
rect 172348 68814 172376 71726
rect 173084 69154 173112 71726
rect 173072 69148 173124 69154
rect 173072 69090 173124 69096
rect 173164 69080 173216 69086
rect 173164 69022 173216 69028
rect 172336 68808 172388 68814
rect 172336 68750 172388 68756
rect 173176 16046 173204 69022
rect 173256 16108 173308 16114
rect 173256 16050 173308 16056
rect 173164 16040 173216 16046
rect 173164 15982 173216 15988
rect 171048 12232 171100 12238
rect 171048 12174 171100 12180
rect 171968 4548 172020 4554
rect 171968 4490 172020 4496
rect 170772 3868 170824 3874
rect 170772 3810 170824 3816
rect 170404 3188 170456 3194
rect 170404 3130 170456 3136
rect 170784 480 170812 3810
rect 171980 480 172008 4490
rect 173268 3806 173296 16050
rect 173624 13728 173676 13734
rect 173624 13670 173676 13676
rect 173256 3800 173308 3806
rect 173256 3742 173308 3748
rect 173636 3398 173664 13670
rect 173728 13394 173756 71726
rect 173808 69148 173860 69154
rect 173808 69090 173860 69096
rect 173820 13462 173848 69090
rect 174464 69086 174492 71726
rect 174452 69080 174504 69086
rect 174452 69022 174504 69028
rect 175096 69080 175148 69086
rect 175096 69022 175148 69028
rect 175108 47598 175136 69022
rect 175096 47592 175148 47598
rect 175096 47534 175148 47540
rect 175096 17264 175148 17270
rect 175096 17206 175148 17212
rect 173808 13456 173860 13462
rect 173808 13398 173860 13404
rect 173716 13388 173768 13394
rect 173716 13330 173768 13336
rect 175108 3398 175136 17206
rect 175200 14686 175228 71726
rect 175844 69086 175872 71726
rect 175832 69080 175884 69086
rect 175832 69022 175884 69028
rect 176476 69080 176528 69086
rect 176476 69022 176528 69028
rect 176488 49026 176516 69022
rect 176476 49020 176528 49026
rect 176476 48962 176528 48968
rect 175188 14680 175240 14686
rect 175188 14622 175240 14628
rect 176580 11966 176608 71726
rect 177224 68746 177252 71726
rect 177776 71726 177942 71754
rect 178604 71726 178640 71754
rect 179310 71754 179338 72012
rect 180008 71754 180036 72012
rect 179310 71726 179368 71754
rect 177212 68740 177264 68746
rect 177212 68682 177264 68688
rect 177304 68604 177356 68610
rect 177304 68546 177356 68552
rect 176568 11960 176620 11966
rect 176568 11902 176620 11908
rect 175464 4616 175516 4622
rect 175464 4558 175516 4564
rect 173164 3392 173216 3398
rect 173164 3334 173216 3340
rect 173624 3392 173676 3398
rect 173624 3334 173676 3340
rect 174268 3392 174320 3398
rect 174268 3334 174320 3340
rect 175096 3392 175148 3398
rect 175096 3334 175148 3340
rect 173176 480 173204 3334
rect 174280 480 174308 3334
rect 175476 480 175504 4558
rect 177316 3942 177344 68546
rect 177776 13326 177804 71726
rect 178604 69086 178632 71726
rect 178592 69080 178644 69086
rect 178592 69022 178644 69028
rect 179236 69080 179288 69086
rect 179236 69022 179288 69028
rect 177856 17468 177908 17474
rect 177856 17410 177908 17416
rect 177764 13320 177816 13326
rect 177764 13262 177816 13268
rect 177304 3936 177356 3942
rect 177304 3878 177356 3884
rect 177868 3398 177896 17410
rect 178684 17332 178736 17338
rect 178684 17274 178736 17280
rect 178696 3874 178724 17274
rect 179248 14618 179276 69022
rect 179236 14612 179288 14618
rect 179236 14554 179288 14560
rect 179340 7070 179368 71726
rect 179984 71726 180036 71754
rect 180705 71754 180733 72012
rect 181403 71754 181431 72012
rect 182101 71754 182129 72012
rect 180705 71726 180748 71754
rect 181403 71726 181484 71754
rect 179984 69086 180012 71726
rect 179972 69080 180024 69086
rect 179972 69022 180024 69028
rect 180616 69080 180668 69086
rect 180616 69022 180668 69028
rect 180248 9512 180300 9518
rect 180248 9454 180300 9460
rect 179328 7064 179380 7070
rect 179328 7006 179380 7012
rect 179052 4684 179104 4690
rect 179052 4626 179104 4632
rect 178684 3868 178736 3874
rect 178684 3810 178736 3816
rect 177948 3800 178000 3806
rect 177948 3742 178000 3748
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 177856 3392 177908 3398
rect 177856 3334 177908 3340
rect 176672 480 176700 3334
rect 177960 1986 177988 3742
rect 177868 1958 177988 1986
rect 177868 480 177896 1958
rect 179064 480 179092 4626
rect 180260 480 180288 9454
rect 180628 7138 180656 69022
rect 180720 7206 180748 71726
rect 181456 69086 181484 71726
rect 182008 71726 182129 71754
rect 182799 71754 182827 72012
rect 183497 71754 183525 72012
rect 182799 71726 182864 71754
rect 181444 69080 181496 69086
rect 181444 69022 181496 69028
rect 181904 12368 181956 12374
rect 181904 12310 181956 12316
rect 180708 7200 180760 7206
rect 180708 7142 180760 7148
rect 180616 7132 180668 7138
rect 180616 7074 180668 7080
rect 181916 3398 181944 12310
rect 182008 7342 182036 71726
rect 182836 69086 182864 71726
rect 183480 71726 183525 71754
rect 184194 71754 184222 72012
rect 184892 71754 184920 72012
rect 184194 71726 184244 71754
rect 182088 69080 182140 69086
rect 182088 69022 182140 69028
rect 182824 69080 182876 69086
rect 182824 69022 182876 69028
rect 183376 69080 183428 69086
rect 183376 69022 183428 69028
rect 181996 7336 182048 7342
rect 181996 7278 182048 7284
rect 182100 7274 182128 69022
rect 183388 7410 183416 69022
rect 183480 7478 183508 71726
rect 184216 69086 184244 71726
rect 184768 71726 184920 71754
rect 185590 71754 185618 72012
rect 186288 71754 186316 72012
rect 186986 71754 187014 72012
rect 185590 71726 185624 71754
rect 186288 71726 186360 71754
rect 184204 69080 184256 69086
rect 184204 69022 184256 69028
rect 183744 9308 183796 9314
rect 183744 9250 183796 9256
rect 183468 7472 183520 7478
rect 183468 7414 183520 7420
rect 183376 7404 183428 7410
rect 183376 7346 183428 7352
rect 182088 7268 182140 7274
rect 182088 7210 182140 7216
rect 182548 4752 182600 4758
rect 182548 4694 182600 4700
rect 181444 3392 181496 3398
rect 181444 3334 181496 3340
rect 181904 3392 181956 3398
rect 181904 3334 181956 3340
rect 181456 480 181484 3334
rect 182560 480 182588 4694
rect 183756 480 183784 9250
rect 184768 8294 184796 71726
rect 185596 69086 185624 71726
rect 186332 69154 186360 71726
rect 186976 71726 187014 71754
rect 187683 71754 187711 72012
rect 188381 71754 188409 72012
rect 187683 71726 187740 71754
rect 186320 69148 186372 69154
rect 186320 69090 186372 69096
rect 186976 69086 187004 71726
rect 187712 69154 187740 71726
rect 188356 71726 188409 71754
rect 189079 71754 189107 72012
rect 189777 71754 189805 72012
rect 190475 71754 190503 72012
rect 189079 71726 189120 71754
rect 189777 71726 189856 71754
rect 187608 69148 187660 69154
rect 187608 69090 187660 69096
rect 187700 69148 187752 69154
rect 187700 69090 187752 69096
rect 184848 69080 184900 69086
rect 184848 69022 184900 69028
rect 185584 69080 185636 69086
rect 185584 69022 185636 69028
rect 186228 69080 186280 69086
rect 186228 69022 186280 69028
rect 186964 69080 187016 69086
rect 186964 69022 187016 69028
rect 187516 69080 187568 69086
rect 187516 69022 187568 69028
rect 184756 8288 184808 8294
rect 184756 8230 184808 8236
rect 184860 7546 184888 69022
rect 186240 8226 186268 69022
rect 187332 10804 187384 10810
rect 187332 10746 187384 10752
rect 186228 8220 186280 8226
rect 186228 8162 186280 8168
rect 184848 7540 184900 7546
rect 184848 7482 184900 7488
rect 186136 5500 186188 5506
rect 186136 5442 186188 5448
rect 184940 3868 184992 3874
rect 184940 3810 184992 3816
rect 184952 480 184980 3810
rect 186148 480 186176 5442
rect 187344 480 187372 10746
rect 187528 8090 187556 69022
rect 187620 8158 187648 69090
rect 188356 69086 188384 71726
rect 189092 69154 189120 71726
rect 188896 69148 188948 69154
rect 188896 69090 188948 69096
rect 189080 69148 189132 69154
rect 189080 69090 189132 69096
rect 188344 69080 188396 69086
rect 188344 69022 188396 69028
rect 187608 8152 187660 8158
rect 187608 8094 187660 8100
rect 187516 8084 187568 8090
rect 187516 8026 187568 8032
rect 188908 8022 188936 69090
rect 189828 69086 189856 71726
rect 190472 71726 190503 71754
rect 191172 71754 191200 72012
rect 191870 71754 191898 72012
rect 191172 71726 191236 71754
rect 190472 69154 190500 71726
rect 190276 69148 190328 69154
rect 190276 69090 190328 69096
rect 190460 69148 190512 69154
rect 190460 69090 190512 69096
rect 188988 69080 189040 69086
rect 188988 69022 189040 69028
rect 189816 69080 189868 69086
rect 189816 69022 189868 69028
rect 188896 8016 188948 8022
rect 188896 7958 188948 7964
rect 189000 7954 189028 69022
rect 188988 7948 189040 7954
rect 188988 7890 189040 7896
rect 190288 7886 190316 69090
rect 191208 69086 191236 71726
rect 191852 71726 191898 71754
rect 192568 71754 192596 72012
rect 193266 71754 193294 72012
rect 193964 71754 193992 72012
rect 194661 71754 194689 72012
rect 195359 71754 195387 72012
rect 192568 71726 192616 71754
rect 193266 71726 193352 71754
rect 193964 71726 193996 71754
rect 194661 71726 194732 71754
rect 191656 69148 191708 69154
rect 191656 69090 191708 69096
rect 190368 69080 190420 69086
rect 190368 69022 190420 69028
rect 191196 69080 191248 69086
rect 191196 69022 191248 69028
rect 190276 7880 190328 7886
rect 190276 7822 190328 7828
rect 190380 7818 190408 69022
rect 191564 10872 191616 10878
rect 191564 10814 191616 10820
rect 190368 7812 190420 7818
rect 190368 7754 190420 7760
rect 189724 5432 189776 5438
rect 189724 5374 189776 5380
rect 188528 4004 188580 4010
rect 188528 3946 188580 3952
rect 188540 480 188568 3946
rect 189736 480 189764 5374
rect 191576 2922 191604 10814
rect 191668 7750 191696 69090
rect 191852 69086 191880 71726
rect 191748 69080 191800 69086
rect 191748 69022 191800 69028
rect 191840 69080 191892 69086
rect 191840 69022 191892 69028
rect 191656 7744 191708 7750
rect 191656 7686 191708 7692
rect 191760 7682 191788 69022
rect 192588 67046 192616 71726
rect 193324 69698 193352 71726
rect 193312 69692 193364 69698
rect 193312 69634 193364 69640
rect 193128 69080 193180 69086
rect 193128 69022 193180 69028
rect 192576 67040 192628 67046
rect 192576 66982 192628 66988
rect 191748 7676 191800 7682
rect 191748 7618 191800 7624
rect 193140 7614 193168 69022
rect 193968 68542 193996 71726
rect 194704 69154 194732 71726
rect 195348 71726 195387 71754
rect 196057 71754 196085 72012
rect 196755 71754 196783 72012
rect 196057 71726 196112 71754
rect 194692 69148 194744 69154
rect 194692 69090 194744 69096
rect 195348 69086 195376 71726
rect 196084 69154 196112 71726
rect 196728 71726 196783 71754
rect 197453 71754 197481 72012
rect 198150 71754 198178 72012
rect 198848 71754 198876 72012
rect 197453 71726 197492 71754
rect 198150 71726 198228 71754
rect 195888 69148 195940 69154
rect 195888 69090 195940 69096
rect 196072 69148 196124 69154
rect 196072 69090 196124 69096
rect 195336 69080 195388 69086
rect 195336 69022 195388 69028
rect 195796 69080 195848 69086
rect 195796 69022 195848 69028
rect 193956 68536 194008 68542
rect 193956 68478 194008 68484
rect 195244 17400 195296 17406
rect 195244 17342 195296 17348
rect 193128 7608 193180 7614
rect 193128 7550 193180 7556
rect 193220 5364 193272 5370
rect 193220 5306 193272 5312
rect 192024 3936 192076 3942
rect 192024 3878 192076 3884
rect 190828 2916 190880 2922
rect 190828 2858 190880 2864
rect 191564 2916 191616 2922
rect 191564 2858 191616 2864
rect 190840 480 190868 2858
rect 192036 480 192064 3878
rect 193232 480 193260 5306
rect 194416 4208 194468 4214
rect 194416 4150 194468 4156
rect 194428 480 194456 4150
rect 195256 4010 195284 17342
rect 195336 14816 195388 14822
rect 195336 14758 195388 14764
rect 195244 4004 195296 4010
rect 195244 3946 195296 3952
rect 195348 3806 195376 14758
rect 195808 14482 195836 69022
rect 195796 14476 195848 14482
rect 195796 14418 195848 14424
rect 195612 13660 195664 13666
rect 195612 13602 195664 13608
rect 195336 3800 195388 3806
rect 195336 3742 195388 3748
rect 195624 480 195652 13602
rect 195900 13258 195928 69090
rect 196728 69086 196756 71726
rect 197176 69148 197228 69154
rect 197176 69090 197228 69096
rect 196716 69080 196768 69086
rect 196716 69022 196768 69028
rect 196624 16176 196676 16182
rect 196624 16118 196676 16124
rect 195888 13252 195940 13258
rect 195888 13194 195940 13200
rect 196636 3874 196664 16118
rect 197188 15910 197216 69090
rect 197268 69080 197320 69086
rect 197268 69022 197320 69028
rect 197176 15904 197228 15910
rect 197176 15846 197228 15852
rect 197280 11830 197308 69022
rect 197464 65618 197492 71726
rect 198004 69216 198056 69222
rect 198004 69158 198056 69164
rect 197452 65612 197504 65618
rect 197452 65554 197504 65560
rect 197268 11824 197320 11830
rect 197268 11766 197320 11772
rect 196808 5296 196860 5302
rect 196808 5238 196860 5244
rect 196624 3868 196676 3874
rect 196624 3810 196676 3816
rect 196820 480 196848 5238
rect 198016 4214 198044 69158
rect 198200 69086 198228 71726
rect 198844 71726 198876 71754
rect 199546 71754 199574 72012
rect 200244 71754 200272 72012
rect 199546 71726 199608 71754
rect 198844 69154 198872 71726
rect 198832 69148 198884 69154
rect 198832 69090 198884 69096
rect 199580 69086 199608 71726
rect 200224 71726 200272 71754
rect 200942 71754 200970 72012
rect 201639 71754 201667 72012
rect 202337 71754 202365 72012
rect 203035 71754 203063 72012
rect 203733 71754 203761 72012
rect 200942 71726 201356 71754
rect 201639 71726 201724 71754
rect 202337 71726 202736 71754
rect 203035 71726 203104 71754
rect 199936 69148 199988 69154
rect 199936 69090 199988 69096
rect 198188 69080 198240 69086
rect 198188 69022 198240 69028
rect 198648 69080 198700 69086
rect 198648 69022 198700 69028
rect 199568 69080 199620 69086
rect 199568 69022 199620 69028
rect 198556 18828 198608 18834
rect 198556 18770 198608 18776
rect 198004 4208 198056 4214
rect 198004 4150 198056 4156
rect 198568 3398 198596 18770
rect 198660 13190 198688 69022
rect 198648 13184 198700 13190
rect 198648 13126 198700 13132
rect 199948 9586 199976 69090
rect 200224 69086 200252 71726
rect 200028 69080 200080 69086
rect 200028 69022 200080 69028
rect 200212 69080 200264 69086
rect 200212 69022 200264 69028
rect 199936 9580 199988 9586
rect 199936 9522 199988 9528
rect 200040 9450 200068 69022
rect 200028 9444 200080 9450
rect 200028 9386 200080 9392
rect 201328 9178 201356 71726
rect 201696 69086 201724 71726
rect 201408 69080 201460 69086
rect 201408 69022 201460 69028
rect 201684 69080 201736 69086
rect 201684 69022 201736 69028
rect 201420 9382 201448 69022
rect 202604 18692 202656 18698
rect 202604 18634 202656 18640
rect 202512 10940 202564 10946
rect 202512 10882 202564 10888
rect 201408 9376 201460 9382
rect 201408 9318 201460 9324
rect 201316 9172 201368 9178
rect 201316 9114 201368 9120
rect 200304 5228 200356 5234
rect 200304 5170 200356 5176
rect 199108 3800 199160 3806
rect 199108 3742 199160 3748
rect 197912 3392 197964 3398
rect 197912 3334 197964 3340
rect 198556 3392 198608 3398
rect 198556 3334 198608 3340
rect 197924 480 197952 3334
rect 199120 480 199148 3742
rect 200316 480 200344 5170
rect 202524 3126 202552 10882
rect 202616 6914 202644 18634
rect 202708 9042 202736 71726
rect 203076 69086 203104 71726
rect 203720 71726 203761 71754
rect 204431 71754 204459 72012
rect 205128 71754 205156 72012
rect 204431 71726 204484 71754
rect 203720 69154 203748 71726
rect 203708 69148 203760 69154
rect 203708 69090 203760 69096
rect 202788 69080 202840 69086
rect 202788 69022 202840 69028
rect 203064 69080 203116 69086
rect 203064 69022 203116 69028
rect 204168 69080 204220 69086
rect 204168 69022 204220 69028
rect 202800 9110 202828 69022
rect 202788 9104 202840 9110
rect 202788 9046 202840 9052
rect 202696 9036 202748 9042
rect 202696 8978 202748 8984
rect 204180 8974 204208 69022
rect 204456 68474 204484 71726
rect 205100 71726 205156 71754
rect 205826 71754 205854 72012
rect 206524 71754 206552 72012
rect 207222 71754 207250 72012
rect 205826 71726 205864 71754
rect 206524 71726 206968 71754
rect 204996 69828 205048 69834
rect 204996 69770 205048 69776
rect 204904 69352 204956 69358
rect 204904 69294 204956 69300
rect 204444 68468 204496 68474
rect 204444 68410 204496 68416
rect 204168 8968 204220 8974
rect 204168 8910 204220 8916
rect 202616 6886 202736 6914
rect 201500 3120 201552 3126
rect 201500 3062 201552 3068
rect 202512 3120 202564 3126
rect 202512 3062 202564 3068
rect 201512 480 201540 3062
rect 202708 480 202736 6886
rect 204916 6730 204944 69294
rect 204904 6724 204956 6730
rect 204904 6666 204956 6672
rect 205008 6118 205036 69770
rect 205100 69698 205128 71726
rect 205088 69692 205140 69698
rect 205088 69634 205140 69640
rect 205836 66978 205864 71726
rect 206284 69420 206336 69426
rect 206284 69362 206336 69368
rect 205824 66972 205876 66978
rect 205824 66914 205876 66920
rect 206296 6866 206324 69362
rect 206376 14884 206428 14890
rect 206376 14826 206428 14832
rect 206284 6860 206336 6866
rect 206284 6802 206336 6808
rect 205088 6792 205140 6798
rect 205088 6734 205140 6740
rect 204996 6112 205048 6118
rect 204996 6054 205048 6060
rect 203892 5160 203944 5166
rect 203892 5102 203944 5108
rect 203904 480 203932 5102
rect 205100 480 205128 6734
rect 206388 3942 206416 14826
rect 206940 13122 206968 71726
rect 207216 71726 207250 71754
rect 207920 71754 207948 72012
rect 208617 71754 208645 72012
rect 207920 71726 207980 71754
rect 207216 69358 207244 71726
rect 207204 69352 207256 69358
rect 207204 69294 207256 69300
rect 207952 69154 207980 71726
rect 208596 71726 208645 71754
rect 209315 71754 209343 72012
rect 210013 71754 210041 72012
rect 210711 71754 210739 72012
rect 211409 71754 211437 72012
rect 212106 71754 212134 72012
rect 212804 71754 212832 72012
rect 213502 71754 213530 72012
rect 214200 71754 214228 72012
rect 214898 71754 214926 72012
rect 215595 71754 215623 72012
rect 209315 71726 209360 71754
rect 210013 71726 210096 71754
rect 210711 71726 211108 71754
rect 211409 71726 211476 71754
rect 212106 71726 212488 71754
rect 212804 71726 212856 71754
rect 213502 71726 213776 71754
rect 214200 71726 214236 71754
rect 214898 71726 215248 71754
rect 208596 69834 208624 71726
rect 208584 69828 208636 69834
rect 208584 69770 208636 69776
rect 209136 69284 209188 69290
rect 209136 69226 209188 69232
rect 207940 69148 207992 69154
rect 207940 69090 207992 69096
rect 209044 67244 209096 67250
rect 209044 67186 209096 67192
rect 206928 13116 206980 13122
rect 206928 13058 206980 13064
rect 207388 5092 207440 5098
rect 207388 5034 207440 5040
rect 206376 3936 206428 3942
rect 206376 3878 206428 3884
rect 206192 3868 206244 3874
rect 206192 3810 206244 3816
rect 206204 480 206232 3810
rect 207400 480 207428 5034
rect 209056 3806 209084 67186
rect 209148 10742 209176 69226
rect 209332 66910 209360 71726
rect 209688 69420 209740 69426
rect 209688 69362 209740 69368
rect 209320 66904 209372 66910
rect 209320 66846 209372 66852
rect 209136 10736 209188 10742
rect 209136 10678 209188 10684
rect 209044 3800 209096 3806
rect 209044 3742 209096 3748
rect 209700 3398 209728 69362
rect 210068 69086 210096 71726
rect 210056 69080 210108 69086
rect 210056 69022 210108 69028
rect 210976 69080 211028 69086
rect 210976 69022 211028 69028
rect 210988 6914 211016 69022
rect 210896 6886 211016 6914
rect 210896 4350 210924 6886
rect 210976 5024 211028 5030
rect 210976 4966 211028 4972
rect 210884 4344 210936 4350
rect 210884 4286 210936 4292
rect 209780 3936 209832 3942
rect 209780 3878 209832 3884
rect 208584 3392 208636 3398
rect 208584 3334 208636 3340
rect 209688 3392 209740 3398
rect 209688 3334 209740 3340
rect 208596 480 208624 3334
rect 209792 480 209820 3878
rect 210988 480 211016 4966
rect 211080 4418 211108 71726
rect 211448 69086 211476 71726
rect 211436 69080 211488 69086
rect 211436 69022 211488 69028
rect 212356 69080 212408 69086
rect 212356 69022 212408 69028
rect 212172 5908 212224 5914
rect 212172 5850 212224 5856
rect 211068 4412 211120 4418
rect 211068 4354 211120 4360
rect 212184 480 212212 5850
rect 212368 4486 212396 69022
rect 212460 4554 212488 71726
rect 212828 69086 212856 71726
rect 213552 69148 213604 69154
rect 213552 69090 213604 69096
rect 212816 69080 212868 69086
rect 212816 69022 212868 69028
rect 213564 68406 213592 69090
rect 213552 68400 213604 68406
rect 213552 68342 213604 68348
rect 213748 4690 213776 71726
rect 214208 69086 214236 71726
rect 213828 69080 213880 69086
rect 213828 69022 213880 69028
rect 214196 69080 214248 69086
rect 214196 69022 214248 69028
rect 215116 69080 215168 69086
rect 215116 69022 215168 69028
rect 213736 4684 213788 4690
rect 213736 4626 213788 4632
rect 213840 4622 213868 69022
rect 214472 4956 214524 4962
rect 214472 4898 214524 4904
rect 213828 4616 213880 4622
rect 213828 4558 213880 4564
rect 212448 4548 212500 4554
rect 212448 4490 212500 4496
rect 212356 4480 212408 4486
rect 212356 4422 212408 4428
rect 213368 3800 213420 3806
rect 213368 3742 213420 3748
rect 213380 480 213408 3742
rect 214484 480 214512 4898
rect 215128 4758 215156 69022
rect 215220 5506 215248 71726
rect 215588 71726 215623 71754
rect 216293 71754 216321 72012
rect 216991 71754 217019 72012
rect 216293 71726 216628 71754
rect 215588 69086 215616 71726
rect 215576 69080 215628 69086
rect 215576 69022 215628 69028
rect 216496 69080 216548 69086
rect 216496 69022 216548 69028
rect 215668 9648 215720 9654
rect 215668 9590 215720 9596
rect 215208 5500 215260 5506
rect 215208 5442 215260 5448
rect 215116 4752 215168 4758
rect 215116 4694 215168 4700
rect 215680 480 215708 9590
rect 216508 5438 216536 69022
rect 216496 5432 216548 5438
rect 216496 5374 216548 5380
rect 216600 5370 216628 71726
rect 216968 71726 217019 71754
rect 217689 71754 217717 72012
rect 218387 71754 218415 72012
rect 217689 71726 218008 71754
rect 218387 71726 218468 71754
rect 216968 69086 216996 71726
rect 216956 69080 217008 69086
rect 216956 69022 217008 69028
rect 217876 69080 217928 69086
rect 217876 69022 217928 69028
rect 216588 5364 216640 5370
rect 216588 5306 216640 5312
rect 217888 5302 217916 69022
rect 217876 5296 217928 5302
rect 217876 5238 217928 5244
rect 217980 5234 218008 71726
rect 218440 69086 218468 71726
rect 218428 69080 218480 69086
rect 218428 69022 218480 69028
rect 218980 69080 219032 69086
rect 218980 69022 219032 69028
rect 218992 64874 219020 69022
rect 219084 68490 219112 72012
rect 219782 71754 219810 72012
rect 220480 71754 220508 72012
rect 221178 71754 221206 72012
rect 221876 71754 221904 72012
rect 222573 71890 222601 72012
rect 222573 71862 222608 71890
rect 219782 71726 219848 71754
rect 220480 71726 220768 71754
rect 221178 71726 221228 71754
rect 221876 71726 222056 71754
rect 219820 69086 219848 71726
rect 219808 69080 219860 69086
rect 219808 69022 219860 69028
rect 220636 69080 220688 69086
rect 220636 69022 220688 69028
rect 219084 68462 219388 68490
rect 218992 64846 219296 64874
rect 219268 6914 219296 64846
rect 219176 6886 219296 6914
rect 217968 5228 218020 5234
rect 217968 5170 218020 5176
rect 219176 5166 219204 6886
rect 219256 5976 219308 5982
rect 219256 5918 219308 5924
rect 219164 5160 219216 5166
rect 219164 5102 219216 5108
rect 218060 4888 218112 4894
rect 218060 4830 218112 4836
rect 216864 4072 216916 4078
rect 216864 4014 216916 4020
rect 216876 480 216904 4014
rect 218072 480 218100 4830
rect 219268 480 219296 5918
rect 219360 5098 219388 68462
rect 219348 5092 219400 5098
rect 219348 5034 219400 5040
rect 220648 5030 220676 69022
rect 220636 5024 220688 5030
rect 220636 4966 220688 4972
rect 220740 4962 220768 71726
rect 221200 69086 221228 71726
rect 221188 69080 221240 69086
rect 221188 69022 221240 69028
rect 220728 4956 220780 4962
rect 220728 4898 220780 4904
rect 222028 4826 222056 71726
rect 222108 69080 222160 69086
rect 222108 69022 222160 69028
rect 222120 4894 222148 69022
rect 222580 65550 222608 71862
rect 223271 71754 223299 72012
rect 223969 71754 223997 72012
rect 222764 71726 223299 71754
rect 223960 71726 223997 71754
rect 224667 71754 224695 72012
rect 225365 71754 225393 72012
rect 224667 71726 224724 71754
rect 222568 65544 222620 65550
rect 222568 65486 222620 65492
rect 222764 64874 222792 71726
rect 223960 69902 223988 71726
rect 224696 70038 224724 71726
rect 225340 71726 225393 71754
rect 226062 71754 226090 72012
rect 226760 71754 226788 72012
rect 227458 71754 227486 72012
rect 228156 71754 228184 72012
rect 228854 71754 228882 72012
rect 226062 71726 226104 71754
rect 225340 70174 225368 71726
rect 226076 70310 226104 71726
rect 226720 71726 226788 71754
rect 227456 71726 227486 71754
rect 227824 71726 228184 71754
rect 228836 71726 228882 71754
rect 229551 71754 229579 72012
rect 230249 71754 230277 72012
rect 229551 71726 229600 71754
rect 226064 70304 226116 70310
rect 226064 70246 226116 70252
rect 226720 70242 226748 71726
rect 227456 70378 227484 71726
rect 227444 70372 227496 70378
rect 227444 70314 227496 70320
rect 226708 70236 226760 70242
rect 226708 70178 226760 70184
rect 225328 70168 225380 70174
rect 225328 70110 225380 70116
rect 224684 70032 224736 70038
rect 224684 69974 224736 69980
rect 223948 69896 224000 69902
rect 223948 69838 224000 69844
rect 227628 69624 227680 69630
rect 227628 69566 227680 69572
rect 224224 69556 224276 69562
rect 224224 69498 224276 69504
rect 222844 69284 222896 69290
rect 222844 69226 222896 69232
rect 222212 64846 222792 64874
rect 222212 9246 222240 64846
rect 222856 9518 222884 69226
rect 222936 18760 222988 18766
rect 222936 18702 222988 18708
rect 222844 9512 222896 9518
rect 222844 9454 222896 9460
rect 222200 9240 222252 9246
rect 222200 9182 222252 9188
rect 222752 9240 222804 9246
rect 222752 9182 222804 9188
rect 222108 4888 222160 4894
rect 222108 4830 222160 4836
rect 221556 4820 221608 4826
rect 221556 4762 221608 4768
rect 222016 4820 222068 4826
rect 222016 4762 222068 4768
rect 220452 2916 220504 2922
rect 220452 2858 220504 2864
rect 220464 480 220492 2858
rect 221568 480 221596 4762
rect 222764 480 222792 9182
rect 222948 2922 222976 18702
rect 224236 6050 224264 69498
rect 226984 69488 227036 69494
rect 226984 69430 227036 69436
rect 224316 69352 224368 69358
rect 224316 69294 224368 69300
rect 224328 11762 224356 69294
rect 224408 16244 224460 16250
rect 224408 16186 224460 16192
rect 224316 11756 224368 11762
rect 224316 11698 224368 11704
rect 224224 6044 224276 6050
rect 224224 5986 224276 5992
rect 223948 4004 224000 4010
rect 223948 3946 224000 3952
rect 222936 2916 222988 2922
rect 222936 2858 222988 2864
rect 223960 480 223988 3946
rect 224420 3874 224448 16186
rect 226996 11694 227024 69430
rect 227076 22772 227128 22778
rect 227076 22714 227128 22720
rect 226984 11688 227036 11694
rect 226984 11630 227036 11636
rect 225144 4276 225196 4282
rect 225144 4218 225196 4224
rect 224408 3868 224460 3874
rect 224408 3810 224460 3816
rect 225156 480 225184 4218
rect 227088 4078 227116 22714
rect 227076 4072 227128 4078
rect 227076 4014 227128 4020
rect 227536 3936 227588 3942
rect 227536 3878 227588 3884
rect 226340 3392 226392 3398
rect 226340 3334 226392 3340
rect 226352 480 226380 3334
rect 227548 480 227576 3878
rect 227640 3398 227668 69566
rect 227824 12102 227852 71726
rect 228364 69896 228416 69902
rect 228364 69838 228416 69844
rect 227812 12096 227864 12102
rect 227812 12038 227864 12044
rect 228376 10674 228404 69838
rect 228836 69562 228864 71726
rect 228824 69556 228876 69562
rect 228824 69498 228876 69504
rect 229572 68610 229600 71726
rect 230216 71726 230277 71754
rect 230480 71800 230532 71806
rect 230947 71754 230975 72012
rect 231645 71806 231673 72012
rect 230480 71742 230532 71748
rect 230216 69902 230244 71726
rect 230204 69896 230256 69902
rect 230204 69838 230256 69844
rect 229560 68604 229612 68610
rect 229560 68546 229612 68552
rect 228456 44872 228508 44878
rect 228456 44814 228508 44820
rect 228364 10668 228416 10674
rect 228364 10610 228416 10616
rect 228468 3874 228496 44814
rect 230492 12170 230520 71742
rect 230584 71726 230975 71754
rect 231633 71800 231685 71806
rect 232343 71754 232371 72012
rect 233040 71754 233068 72012
rect 233738 71890 233766 72012
rect 231633 71742 231685 71748
rect 231872 71726 232371 71754
rect 232424 71726 233068 71754
rect 233252 71862 233766 71890
rect 230584 14550 230612 71726
rect 231124 70168 231176 70174
rect 231124 70110 231176 70116
rect 230572 14544 230624 14550
rect 230572 14486 230624 14492
rect 230480 12164 230532 12170
rect 230480 12106 230532 12112
rect 228732 6112 228784 6118
rect 228732 6054 228784 6060
rect 229836 6112 229888 6118
rect 229836 6054 229888 6060
rect 228456 3868 228508 3874
rect 228456 3810 228508 3816
rect 227628 3392 227680 3398
rect 227628 3334 227680 3340
rect 228744 480 228772 6054
rect 229848 480 229876 6054
rect 231136 5914 231164 70110
rect 231216 14952 231268 14958
rect 231216 14894 231268 14900
rect 231124 5908 231176 5914
rect 231124 5850 231176 5856
rect 231228 3942 231256 14894
rect 231872 13734 231900 71726
rect 232424 64874 232452 71726
rect 233252 69290 233280 71862
rect 234436 71754 234464 72012
rect 233344 71726 234464 71754
rect 234712 71800 234764 71806
rect 235134 71754 235162 72012
rect 235832 71806 235860 72012
rect 234712 71742 234764 71748
rect 233240 69284 233292 69290
rect 233240 69226 233292 69232
rect 232504 69080 232556 69086
rect 232504 69022 232556 69028
rect 231964 64846 232452 64874
rect 231964 17474 231992 64846
rect 231952 17468 232004 17474
rect 231952 17410 232004 17416
rect 231860 13728 231912 13734
rect 231860 13670 231912 13676
rect 231768 13592 231820 13598
rect 231768 13534 231820 13540
rect 231216 3936 231268 3942
rect 231216 3878 231268 3884
rect 231780 3398 231808 13534
rect 232516 10810 232544 69022
rect 232596 17468 232648 17474
rect 232596 17410 232648 17416
rect 232504 10804 232556 10810
rect 232504 10746 232556 10752
rect 232228 6860 232280 6866
rect 232228 6802 232280 6808
rect 231032 3392 231084 3398
rect 231032 3334 231084 3340
rect 231768 3392 231820 3398
rect 231768 3334 231820 3340
rect 231044 480 231072 3334
rect 232240 480 232268 6802
rect 232608 3806 232636 17410
rect 233344 9314 233372 71726
rect 234528 70032 234580 70038
rect 234528 69974 234580 69980
rect 233332 9308 233384 9314
rect 233332 9250 233384 9256
rect 232596 3800 232648 3806
rect 232596 3742 232648 3748
rect 234540 3398 234568 69974
rect 234724 10878 234752 71742
rect 235092 71726 235162 71754
rect 235820 71800 235872 71806
rect 235820 71742 235872 71748
rect 236092 71800 236144 71806
rect 236529 71754 236557 72012
rect 237227 71806 237255 72012
rect 236092 71742 236144 71748
rect 235092 69086 235120 71726
rect 235080 69080 235132 69086
rect 235080 69022 235132 69028
rect 235908 50380 235960 50386
rect 235908 50322 235960 50328
rect 234712 10872 234764 10878
rect 234712 10814 234764 10820
rect 235816 6656 235868 6662
rect 235816 6598 235868 6604
rect 233424 3392 233476 3398
rect 233424 3334 233476 3340
rect 234528 3392 234580 3398
rect 234528 3334 234580 3340
rect 233436 480 233464 3334
rect 234620 3188 234672 3194
rect 234620 3130 234672 3136
rect 234632 480 234660 3130
rect 235828 480 235856 6598
rect 235920 3194 235948 50322
rect 236104 18834 236132 71742
rect 236472 71726 236557 71754
rect 237215 71800 237267 71806
rect 237215 71742 237267 71748
rect 237380 71800 237432 71806
rect 237925 71754 237953 72012
rect 238623 71806 238651 72012
rect 237380 71742 237432 71748
rect 236472 69222 236500 71726
rect 236460 69216 236512 69222
rect 236460 69158 236512 69164
rect 236092 18828 236144 18834
rect 236092 18770 236144 18776
rect 237392 6798 237420 71742
rect 237484 71726 237953 71754
rect 238611 71800 238663 71806
rect 238611 71742 238663 71748
rect 239321 71754 239349 72012
rect 240018 71754 240046 72012
rect 239321 71726 239352 71754
rect 237484 10946 237512 71726
rect 239324 69426 239352 71726
rect 239968 71726 240046 71754
rect 240140 71800 240192 71806
rect 240716 71754 240744 72012
rect 241414 71806 241442 72012
rect 240140 71742 240192 71748
rect 239968 70174 239996 71726
rect 239956 70168 240008 70174
rect 239956 70110 240008 70116
rect 239312 69420 239364 69426
rect 239312 69362 239364 69368
rect 238024 25560 238076 25566
rect 238024 25502 238076 25508
rect 237472 10940 237524 10946
rect 237472 10882 237524 10888
rect 237380 6792 237432 6798
rect 237380 6734 237432 6740
rect 237012 6656 237064 6662
rect 237012 6598 237064 6604
rect 235908 3188 235960 3194
rect 235908 3130 235960 3136
rect 237024 480 237052 6598
rect 238036 4010 238064 25502
rect 239312 6724 239364 6730
rect 239312 6666 239364 6672
rect 238024 4004 238076 4010
rect 238024 3946 238076 3952
rect 238116 3800 238168 3806
rect 238116 3742 238168 3748
rect 238128 480 238156 3742
rect 239324 480 239352 6666
rect 240152 5982 240180 71742
rect 240244 71726 240744 71754
rect 241402 71800 241454 71806
rect 242112 71754 242140 72012
rect 241402 71742 241454 71748
rect 241624 71726 242140 71754
rect 242810 71754 242838 72012
rect 243507 71754 243535 72012
rect 244205 71754 244233 72012
rect 244903 71754 244931 72012
rect 245601 71754 245629 72012
rect 246299 71754 246327 72012
rect 246996 71754 247024 72012
rect 242810 71726 242848 71754
rect 240244 9654 240272 71726
rect 240232 9648 240284 9654
rect 240232 9590 240284 9596
rect 240508 9648 240560 9654
rect 240508 9590 240560 9596
rect 240140 5976 240192 5982
rect 240140 5918 240192 5924
rect 240520 480 240548 9590
rect 241624 9246 241652 71726
rect 242820 69902 242848 71726
rect 243464 71726 243535 71754
rect 244200 71726 244233 71754
rect 244292 71726 244931 71754
rect 245580 71726 245629 71754
rect 245672 71726 246327 71754
rect 246960 71726 247024 71754
rect 247694 71754 247722 72012
rect 248392 71754 248420 72012
rect 249090 71754 249118 72012
rect 247694 71726 247724 71754
rect 248392 71726 248460 71754
rect 242808 69896 242860 69902
rect 242808 69838 242860 69844
rect 243464 69086 243492 71726
rect 244200 70038 244228 71726
rect 244188 70032 244240 70038
rect 244188 69974 244240 69980
rect 242164 69080 242216 69086
rect 242164 69022 242216 69028
rect 243452 69080 243504 69086
rect 243452 69022 243504 69028
rect 241612 9240 241664 9246
rect 241612 9182 241664 9188
rect 242176 6118 242204 69022
rect 242256 17604 242308 17610
rect 242256 17546 242308 17552
rect 242164 6112 242216 6118
rect 242164 6054 242216 6060
rect 242268 3806 242296 17546
rect 244292 6662 244320 71726
rect 245580 68610 245608 71726
rect 244372 68604 244424 68610
rect 244372 68546 244424 68552
rect 245568 68604 245620 68610
rect 245568 68546 245620 68552
rect 244384 9654 244412 68546
rect 244372 9648 244424 9654
rect 244372 9590 244424 9596
rect 244280 6656 244332 6662
rect 244280 6598 244332 6604
rect 242900 6588 242952 6594
rect 242900 6530 242952 6536
rect 242256 3800 242308 3806
rect 242256 3742 242308 3748
rect 241702 3632 241758 3641
rect 241702 3567 241758 3576
rect 241716 480 241744 3567
rect 242912 480 242940 6530
rect 245672 5574 245700 71726
rect 246396 6044 246448 6050
rect 246396 5986 246448 5992
rect 244096 5568 244148 5574
rect 244096 5510 244148 5516
rect 245660 5568 245712 5574
rect 245660 5510 245712 5516
rect 244108 480 244136 5510
rect 245198 3768 245254 3777
rect 245198 3703 245254 3712
rect 245212 480 245240 3703
rect 246408 480 246436 5986
rect 246960 5574 246988 71726
rect 247696 69630 247724 71726
rect 247684 69624 247736 69630
rect 247684 69566 247736 69572
rect 248432 69154 248460 71726
rect 249076 71726 249118 71754
rect 249788 71754 249816 72012
rect 250485 71754 250513 72012
rect 249788 71726 249840 71754
rect 248972 69624 249024 69630
rect 248972 69566 249024 69572
rect 248420 69148 248472 69154
rect 248420 69090 248472 69096
rect 248984 64874 249012 69566
rect 249076 69086 249104 71726
rect 249708 69148 249760 69154
rect 249708 69090 249760 69096
rect 249064 69080 249116 69086
rect 249064 69022 249116 69028
rect 249616 69080 249668 69086
rect 249616 69022 249668 69028
rect 248984 64846 249104 64874
rect 249076 17950 249104 64846
rect 249064 17944 249116 17950
rect 249064 17886 249116 17892
rect 249628 9246 249656 69022
rect 249616 9240 249668 9246
rect 249616 9182 249668 9188
rect 249720 5574 249748 69090
rect 249812 69086 249840 71726
rect 250456 71726 250513 71754
rect 251183 71754 251211 72012
rect 251881 71754 251909 72012
rect 252579 71754 252607 72012
rect 251183 71726 251220 71754
rect 251881 71726 251956 71754
rect 250352 70100 250404 70106
rect 250352 70042 250404 70048
rect 249800 69080 249852 69086
rect 249800 69022 249852 69028
rect 250364 64874 250392 70042
rect 250456 69902 250484 71726
rect 250444 69896 250496 69902
rect 250444 69838 250496 69844
rect 251192 69154 251220 71726
rect 251180 69148 251232 69154
rect 251180 69090 251232 69096
rect 251928 69086 251956 71726
rect 252572 71726 252607 71754
rect 253277 71754 253305 72012
rect 253974 71754 254002 72012
rect 253277 71726 253336 71754
rect 252572 69154 252600 71726
rect 252468 69148 252520 69154
rect 252468 69090 252520 69096
rect 252560 69148 252612 69154
rect 252560 69090 252612 69096
rect 251088 69080 251140 69086
rect 251088 69022 251140 69028
rect 251916 69080 251968 69086
rect 251916 69022 251968 69028
rect 252376 69080 252428 69086
rect 252376 69022 252428 69028
rect 250364 64846 250484 64874
rect 250456 10606 250484 64846
rect 249984 10600 250036 10606
rect 249984 10542 250036 10548
rect 250444 10600 250496 10606
rect 250444 10542 250496 10548
rect 246948 5568 247000 5574
rect 246948 5510 247000 5516
rect 247592 5568 247644 5574
rect 247592 5510 247644 5516
rect 249708 5568 249760 5574
rect 249708 5510 249760 5516
rect 247604 480 247632 5510
rect 248788 3800 248840 3806
rect 248788 3742 248840 3748
rect 248800 480 248828 3742
rect 249996 480 250024 10542
rect 251100 5914 251128 69022
rect 251180 17944 251232 17950
rect 251180 17886 251232 17892
rect 251088 5908 251140 5914
rect 251088 5850 251140 5856
rect 251192 480 251220 17886
rect 252388 5982 252416 69022
rect 252376 5976 252428 5982
rect 252376 5918 252428 5924
rect 252480 4214 252508 69090
rect 253308 69086 253336 71726
rect 253952 71726 254002 71754
rect 254672 71754 254700 72012
rect 255370 71754 255398 72012
rect 254672 71726 254716 71754
rect 255370 71726 255452 71754
rect 253952 69154 253980 71726
rect 253848 69148 253900 69154
rect 253848 69090 253900 69096
rect 253940 69148 253992 69154
rect 253940 69090 253992 69096
rect 253296 69080 253348 69086
rect 253296 69022 253348 69028
rect 253756 69080 253808 69086
rect 253756 69022 253808 69028
rect 253480 10532 253532 10538
rect 253480 10474 253532 10480
rect 252468 4208 252520 4214
rect 252468 4150 252520 4156
rect 252376 3868 252428 3874
rect 252376 3810 252428 3816
rect 252388 480 252416 3810
rect 253492 480 253520 10474
rect 253768 6118 253796 69022
rect 253756 6112 253808 6118
rect 253756 6054 253808 6060
rect 253860 6050 253888 69090
rect 254688 69086 254716 71726
rect 255424 69154 255452 71726
rect 255228 69148 255280 69154
rect 255228 69090 255280 69096
rect 255412 69148 255464 69154
rect 255412 69090 255464 69096
rect 254676 69080 254728 69086
rect 254676 69022 254728 69028
rect 255136 69080 255188 69086
rect 255136 69022 255188 69028
rect 255148 6798 255176 69022
rect 255240 6866 255268 69090
rect 256068 69086 256096 72012
rect 256766 71754 256794 72012
rect 257463 71754 257491 72012
rect 256766 71726 256832 71754
rect 256804 69154 256832 71726
rect 257448 71726 257491 71754
rect 258161 71754 258189 72012
rect 258859 71754 258887 72012
rect 259557 71754 259585 72012
rect 260255 71754 260283 72012
rect 260952 71754 260980 72012
rect 258161 71726 258212 71754
rect 258859 71726 258948 71754
rect 259557 71726 259592 71754
rect 260255 71726 260696 71754
rect 256608 69148 256660 69154
rect 256608 69090 256660 69096
rect 256792 69148 256844 69154
rect 256792 69090 256844 69096
rect 256056 69080 256108 69086
rect 256056 69022 256108 69028
rect 256516 69080 256568 69086
rect 256516 69022 256568 69028
rect 255228 6860 255280 6866
rect 255228 6802 255280 6808
rect 255136 6792 255188 6798
rect 255136 6734 255188 6740
rect 256528 6662 256556 69022
rect 256620 6730 256648 69090
rect 257448 69086 257476 71726
rect 258184 69154 258212 71726
rect 257896 69148 257948 69154
rect 257896 69090 257948 69096
rect 258172 69148 258224 69154
rect 258172 69090 258224 69096
rect 257436 69080 257488 69086
rect 257436 69022 257488 69028
rect 256608 6724 256660 6730
rect 256608 6666 256660 6672
rect 256516 6656 256568 6662
rect 256516 6598 256568 6604
rect 257908 6594 257936 69090
rect 258920 69086 258948 71726
rect 259276 69148 259328 69154
rect 259276 69090 259328 69096
rect 257988 69080 258040 69086
rect 257988 69022 258040 69028
rect 258908 69080 258960 69086
rect 258908 69022 258960 69028
rect 257896 6588 257948 6594
rect 257896 6530 257948 6536
rect 258000 6526 258028 69022
rect 259288 9518 259316 69090
rect 259564 69086 259592 71726
rect 259368 69080 259420 69086
rect 259368 69022 259420 69028
rect 259552 69080 259604 69086
rect 259552 69022 259604 69028
rect 259276 9512 259328 9518
rect 259276 9454 259328 9460
rect 259380 9314 259408 69022
rect 259460 10464 259512 10470
rect 259460 10406 259512 10412
rect 259368 9308 259420 9314
rect 259368 9250 259420 9256
rect 258264 9240 258316 9246
rect 258264 9182 258316 9188
rect 257068 6520 257120 6526
rect 257068 6462 257120 6468
rect 257988 6520 258040 6526
rect 257988 6462 258040 6468
rect 253848 6044 253900 6050
rect 253848 5986 253900 5992
rect 254676 5568 254728 5574
rect 254676 5510 254728 5516
rect 254688 480 254716 5510
rect 255872 3936 255924 3942
rect 255872 3878 255924 3884
rect 255884 480 255912 3878
rect 257080 480 257108 6462
rect 258276 480 258304 9182
rect 259472 3398 259500 10406
rect 260668 8430 260696 71726
rect 260944 71726 260980 71754
rect 261650 71754 261678 72012
rect 262348 71754 262376 72012
rect 261650 71726 261708 71754
rect 260944 69154 260972 71726
rect 260932 69148 260984 69154
rect 260932 69090 260984 69096
rect 261680 69086 261708 71726
rect 262324 71726 262376 71754
rect 263046 71754 263074 72012
rect 263744 71754 263772 72012
rect 264441 71754 264469 72012
rect 265139 71754 265167 72012
rect 265837 71754 265865 72012
rect 263046 71726 263088 71754
rect 263744 71726 263824 71754
rect 264441 71726 264836 71754
rect 265139 71726 265204 71754
rect 262324 69154 262352 71726
rect 262036 69148 262088 69154
rect 262036 69090 262088 69096
rect 262312 69148 262364 69154
rect 262312 69090 262364 69096
rect 260748 69080 260800 69086
rect 260748 69022 260800 69028
rect 261668 69080 261720 69086
rect 261668 69022 261720 69028
rect 260760 9246 260788 69022
rect 260748 9240 260800 9246
rect 260748 9182 260800 9188
rect 262048 8498 262076 69090
rect 263060 69086 263088 71726
rect 263416 69148 263468 69154
rect 263416 69090 263468 69096
rect 262128 69080 262180 69086
rect 262128 69022 262180 69028
rect 263048 69080 263100 69086
rect 263048 69022 263100 69028
rect 262140 8566 262168 69022
rect 263428 8634 263456 69090
rect 263796 69086 263824 71726
rect 263508 69080 263560 69086
rect 263508 69022 263560 69028
rect 263784 69080 263836 69086
rect 263784 69022 263836 69028
rect 263520 8702 263548 69022
rect 264152 10396 264204 10402
rect 264152 10338 264204 10344
rect 263508 8696 263560 8702
rect 263508 8638 263560 8644
rect 263416 8628 263468 8634
rect 263416 8570 263468 8576
rect 262128 8560 262180 8566
rect 262128 8502 262180 8508
rect 262036 8492 262088 8498
rect 262036 8434 262088 8440
rect 260656 8424 260708 8430
rect 260656 8366 260708 8372
rect 261760 5908 261812 5914
rect 261760 5850 261812 5856
rect 259552 4004 259604 4010
rect 259552 3946 259604 3952
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 259564 1986 259592 3946
rect 260656 3392 260708 3398
rect 260656 3334 260708 3340
rect 259472 1958 259592 1986
rect 259472 480 259500 1958
rect 260668 480 260696 3334
rect 261772 480 261800 5850
rect 262956 4072 263008 4078
rect 262956 4014 263008 4020
rect 262968 480 262996 4014
rect 264164 480 264192 10338
rect 264808 8838 264836 71726
rect 264980 69896 265032 69902
rect 264980 69838 265032 69844
rect 264888 69080 264940 69086
rect 264888 69022 264940 69028
rect 264796 8832 264848 8838
rect 264796 8774 264848 8780
rect 264900 8770 264928 69022
rect 264992 16574 265020 69838
rect 265176 69086 265204 71726
rect 265820 71726 265865 71754
rect 266535 71754 266563 72012
rect 267233 71754 267261 72012
rect 267930 71754 267958 72012
rect 268628 71754 268656 72012
rect 269326 71754 269354 72012
rect 266535 71726 266584 71754
rect 267233 71726 267596 71754
rect 267930 71726 267964 71754
rect 268628 71726 268976 71754
rect 265820 70378 265848 71726
rect 265808 70372 265860 70378
rect 265808 70314 265860 70320
rect 266556 69086 266584 71726
rect 265164 69080 265216 69086
rect 265164 69022 265216 69028
rect 266268 69080 266320 69086
rect 266268 69022 266320 69028
rect 266544 69080 266596 69086
rect 266544 69022 266596 69028
rect 264992 16546 265388 16574
rect 264888 8764 264940 8770
rect 264888 8706 264940 8712
rect 265360 480 265388 16546
rect 266280 8906 266308 69022
rect 267568 15026 267596 71726
rect 267936 69086 267964 71726
rect 267648 69080 267700 69086
rect 267648 69022 267700 69028
rect 267924 69080 267976 69086
rect 267924 69022 267976 69028
rect 267556 15020 267608 15026
rect 267556 14962 267608 14968
rect 267660 12442 267688 69022
rect 268948 21418 268976 71726
rect 269316 71726 269354 71754
rect 270024 71754 270052 72012
rect 270722 71754 270750 72012
rect 270024 71726 270448 71754
rect 269316 69086 269344 71726
rect 269028 69080 269080 69086
rect 269028 69022 269080 69028
rect 269304 69080 269356 69086
rect 269304 69022 269356 69028
rect 270316 69080 270368 69086
rect 270316 69022 270368 69028
rect 268936 21412 268988 21418
rect 268936 21354 268988 21360
rect 267648 12436 267700 12442
rect 267648 12378 267700 12384
rect 267740 12028 267792 12034
rect 267740 11970 267792 11976
rect 266268 8900 266320 8906
rect 266268 8842 266320 8848
rect 266544 4140 266596 4146
rect 266544 4082 266596 4088
rect 266556 480 266584 4082
rect 267752 480 267780 11970
rect 269040 4282 269068 69022
rect 270328 16386 270356 69022
rect 270316 16380 270368 16386
rect 270316 16322 270368 16328
rect 270420 13734 270448 71726
rect 270696 71726 270750 71754
rect 271419 71754 271447 72012
rect 272117 71754 272145 72012
rect 272815 71754 272843 72012
rect 273513 71754 273541 72012
rect 274211 71754 274239 72012
rect 274908 71754 274936 72012
rect 275606 71754 275634 72012
rect 276304 71754 276332 72012
rect 277002 71754 277030 72012
rect 277700 71754 277728 72012
rect 271419 71726 271828 71754
rect 272117 71726 272196 71754
rect 272815 71726 273208 71754
rect 273513 71726 273576 71754
rect 274211 71726 274588 71754
rect 274908 71726 274956 71754
rect 275606 71726 275968 71754
rect 276304 71726 276336 71754
rect 277002 71726 277348 71754
rect 270696 69086 270724 71726
rect 270684 69080 270736 69086
rect 270684 69022 270736 69028
rect 271696 69080 271748 69086
rect 271696 69022 271748 69028
rect 271708 17542 271736 69022
rect 271696 17536 271748 17542
rect 271696 17478 271748 17484
rect 271800 16318 271828 71726
rect 272168 69630 272196 71726
rect 272156 69624 272208 69630
rect 272156 69566 272208 69572
rect 271788 16312 271840 16318
rect 271788 16254 271840 16260
rect 270408 13728 270460 13734
rect 270408 13670 270460 13676
rect 271236 10328 271288 10334
rect 271236 10270 271288 10276
rect 268844 4276 268896 4282
rect 268844 4218 268896 4224
rect 269028 4276 269080 4282
rect 269028 4218 269080 4224
rect 268856 480 268884 4218
rect 270040 3392 270092 3398
rect 270040 3334 270092 3340
rect 270052 480 270080 3334
rect 271248 480 271276 10270
rect 273180 9790 273208 71726
rect 273548 69086 273576 71726
rect 274364 69624 274416 69630
rect 274364 69566 274416 69572
rect 273536 69080 273588 69086
rect 273536 69022 273588 69028
rect 274376 67318 274404 69566
rect 274456 69080 274508 69086
rect 274456 69022 274508 69028
rect 274364 67312 274416 67318
rect 274364 67254 274416 67260
rect 274468 9858 274496 69022
rect 274560 9926 274588 71726
rect 274928 69086 274956 71726
rect 274916 69080 274968 69086
rect 274916 69022 274968 69028
rect 275836 69080 275888 69086
rect 275836 69022 275888 69028
rect 274824 10736 274876 10742
rect 274824 10678 274876 10684
rect 274548 9920 274600 9926
rect 274548 9862 274600 9868
rect 274456 9852 274508 9858
rect 274456 9794 274508 9800
rect 273168 9784 273220 9790
rect 273168 9726 273220 9732
rect 272432 5976 272484 5982
rect 272432 5918 272484 5924
rect 272444 480 272472 5918
rect 273628 3324 273680 3330
rect 273628 3266 273680 3272
rect 273640 480 273668 3266
rect 274836 480 274864 10678
rect 275848 9994 275876 69022
rect 275940 10062 275968 71726
rect 276308 69086 276336 71726
rect 276296 69080 276348 69086
rect 276296 69022 276348 69028
rect 277216 69080 277268 69086
rect 277216 69022 277268 69028
rect 277228 10130 277256 69022
rect 277320 10198 277348 71726
rect 277688 71726 277728 71754
rect 278397 71754 278425 72012
rect 279095 71754 279123 72012
rect 278397 71726 278728 71754
rect 277688 69086 277716 71726
rect 277676 69080 277728 69086
rect 277676 69022 277728 69028
rect 278596 69080 278648 69086
rect 278596 69022 278648 69028
rect 278320 10600 278372 10606
rect 278320 10542 278372 10548
rect 277308 10192 277360 10198
rect 277308 10134 277360 10140
rect 277216 10124 277268 10130
rect 277216 10066 277268 10072
rect 275928 10056 275980 10062
rect 275928 9998 275980 10004
rect 275836 9988 275888 9994
rect 275836 9930 275888 9936
rect 276020 6044 276072 6050
rect 276020 5986 276072 5992
rect 276032 480 276060 5986
rect 277124 3256 277176 3262
rect 277124 3198 277176 3204
rect 277136 480 277164 3198
rect 278332 480 278360 10542
rect 278608 10266 278636 69022
rect 278700 11014 278728 71726
rect 279068 71726 279123 71754
rect 279793 71754 279821 72012
rect 280491 71754 280519 72012
rect 281189 71754 281217 72012
rect 281886 71754 281914 72012
rect 282584 71754 282612 72012
rect 283282 71754 283310 72012
rect 283980 71754 284008 72012
rect 284678 71754 284706 72012
rect 285375 71754 285403 72012
rect 286073 71754 286101 72012
rect 279793 71726 280108 71754
rect 280491 71726 280568 71754
rect 281189 71726 281304 71754
rect 281886 71726 281948 71754
rect 282584 71726 282868 71754
rect 283282 71726 283328 71754
rect 283980 71726 284156 71754
rect 284678 71726 284708 71754
rect 285375 71726 285628 71754
rect 279068 69086 279096 71726
rect 279056 69080 279108 69086
rect 279056 69022 279108 69028
rect 279976 69080 280028 69086
rect 279976 69022 280028 69028
rect 278688 11008 278740 11014
rect 278688 10950 278740 10956
rect 279988 10946 280016 69022
rect 279976 10940 280028 10946
rect 279976 10882 280028 10888
rect 280080 10878 280108 71726
rect 280540 69086 280568 71726
rect 280528 69080 280580 69086
rect 280528 69022 280580 69028
rect 280068 10872 280120 10878
rect 280068 10814 280120 10820
rect 281276 10742 281304 71726
rect 281448 70168 281500 70174
rect 281448 70110 281500 70116
rect 281356 69080 281408 69086
rect 281356 69022 281408 69028
rect 281368 10810 281396 69022
rect 281356 10804 281408 10810
rect 281356 10746 281408 10752
rect 281264 10736 281316 10742
rect 281264 10678 281316 10684
rect 278596 10260 278648 10266
rect 278596 10202 278648 10208
rect 279516 6112 279568 6118
rect 279516 6054 279568 6060
rect 279528 480 279556 6054
rect 281460 3126 281488 70110
rect 281920 69086 281948 71726
rect 281908 69080 281960 69086
rect 281908 69022 281960 69028
rect 282736 69080 282788 69086
rect 282736 69022 282788 69028
rect 281908 11688 281960 11694
rect 281908 11630 281960 11636
rect 280712 3120 280764 3126
rect 280712 3062 280764 3068
rect 281448 3120 281500 3126
rect 281448 3062 281500 3068
rect 280724 480 280752 3062
rect 281920 480 281948 11630
rect 282748 10674 282776 69022
rect 282736 10668 282788 10674
rect 282736 10610 282788 10616
rect 282840 10606 282868 71726
rect 283300 69086 283328 71726
rect 283288 69080 283340 69086
rect 283288 69022 283340 69028
rect 282828 10600 282880 10606
rect 282828 10542 282880 10548
rect 284128 10470 284156 71726
rect 284680 69086 284708 71726
rect 284208 69080 284260 69086
rect 284208 69022 284260 69028
rect 284668 69080 284720 69086
rect 284668 69022 284720 69028
rect 285496 69080 285548 69086
rect 285496 69022 285548 69028
rect 284220 10538 284248 69022
rect 285404 11892 285456 11898
rect 285404 11834 285456 11840
rect 284208 10532 284260 10538
rect 284208 10474 284260 10480
rect 284116 10464 284168 10470
rect 284116 10406 284168 10412
rect 283104 6860 283156 6866
rect 283104 6802 283156 6808
rect 283116 480 283144 6802
rect 284300 3188 284352 3194
rect 284300 3130 284352 3136
rect 284312 480 284340 3130
rect 285416 480 285444 11834
rect 285508 10402 285536 69022
rect 285496 10396 285548 10402
rect 285496 10338 285548 10344
rect 285600 10334 285628 71726
rect 286060 71726 286101 71754
rect 286771 71754 286799 72012
rect 287469 71754 287497 72012
rect 286771 71726 287008 71754
rect 286060 69086 286088 71726
rect 286048 69080 286100 69086
rect 286048 69022 286100 69028
rect 286876 69080 286928 69086
rect 286876 69022 286928 69028
rect 286888 12170 286916 69022
rect 286876 12164 286928 12170
rect 286876 12106 286928 12112
rect 286980 12102 287008 71726
rect 287440 71726 287497 71754
rect 288167 71754 288195 72012
rect 288864 71754 288892 72012
rect 289562 71754 289590 72012
rect 288167 71726 288296 71754
rect 288864 71726 288940 71754
rect 287440 69086 287468 71726
rect 287704 70304 287756 70310
rect 287704 70246 287756 70252
rect 287428 69080 287480 69086
rect 287428 69022 287480 69028
rect 287716 13666 287744 70246
rect 288268 64190 288296 71726
rect 288912 69086 288940 71726
rect 289556 71726 289590 71754
rect 290260 71754 290288 72012
rect 290958 71754 290986 72012
rect 290260 71726 290320 71754
rect 289084 69488 289136 69494
rect 289084 69430 289136 69436
rect 288348 69080 288400 69086
rect 288348 69022 288400 69028
rect 288900 69080 288952 69086
rect 288900 69022 288952 69028
rect 288256 64184 288308 64190
rect 288256 64126 288308 64132
rect 287704 13660 287756 13666
rect 287704 13602 287756 13608
rect 286968 12096 287020 12102
rect 286968 12038 287020 12044
rect 288360 12034 288388 69022
rect 288348 12028 288400 12034
rect 288348 11970 288400 11976
rect 285588 10328 285640 10334
rect 285588 10270 285640 10276
rect 286600 6792 286652 6798
rect 286600 6734 286652 6740
rect 286612 480 286640 6734
rect 289096 6458 289124 69430
rect 289556 65754 289584 71726
rect 290292 69358 290320 71726
rect 290936 71726 290986 71754
rect 291656 71754 291684 72012
rect 292353 71754 292381 72012
rect 293051 71754 293079 72012
rect 293749 71754 293777 72012
rect 294447 71754 294475 72012
rect 291656 71726 291700 71754
rect 292353 71726 292528 71754
rect 293051 71726 293080 71754
rect 293749 71726 293816 71754
rect 290280 69352 290332 69358
rect 290280 69294 290332 69300
rect 290936 69086 290964 71726
rect 291672 70242 291700 71726
rect 291660 70236 291712 70242
rect 291660 70178 291712 70184
rect 291844 69556 291896 69562
rect 291844 69498 291896 69504
rect 289728 69080 289780 69086
rect 289728 69022 289780 69028
rect 290924 69080 290976 69086
rect 290924 69022 290976 69028
rect 289544 65748 289596 65754
rect 289544 65690 289596 65696
rect 289740 24138 289768 69022
rect 289728 24132 289780 24138
rect 289728 24074 289780 24080
rect 291856 12374 291884 69498
rect 292396 69352 292448 69358
rect 292396 69294 292448 69300
rect 292408 67114 292436 69294
rect 292396 67108 292448 67114
rect 292396 67050 292448 67056
rect 292500 14550 292528 71726
rect 293052 69426 293080 71726
rect 293788 69630 293816 71726
rect 294432 71726 294475 71754
rect 295145 71754 295173 72012
rect 295842 71754 295870 72012
rect 295145 71726 295196 71754
rect 293776 69624 293828 69630
rect 293776 69566 293828 69572
rect 293040 69420 293092 69426
rect 293040 69362 293092 69368
rect 294432 69290 294460 71726
rect 295168 70038 295196 71726
rect 295812 71726 295870 71754
rect 296540 71754 296568 72012
rect 297238 71754 297266 72012
rect 297936 71754 297964 72012
rect 296540 71726 296668 71754
rect 297238 71726 297312 71754
rect 295812 70106 295840 71726
rect 295984 70372 296036 70378
rect 295984 70314 296036 70320
rect 295800 70100 295852 70106
rect 295800 70042 295852 70048
rect 295156 70032 295208 70038
rect 295156 69974 295208 69980
rect 295248 69352 295300 69358
rect 295248 69294 295300 69300
rect 294420 69284 294472 69290
rect 294420 69226 294472 69232
rect 293776 69080 293828 69086
rect 293776 69022 293828 69028
rect 293788 65686 293816 69022
rect 293776 65680 293828 65686
rect 293776 65622 293828 65628
rect 292488 14544 292540 14550
rect 292488 14486 292540 14492
rect 291844 12368 291896 12374
rect 291844 12310 291896 12316
rect 295260 6914 295288 69294
rect 295892 69284 295944 69290
rect 295892 69226 295944 69232
rect 295904 68610 295932 69226
rect 295892 68604 295944 68610
rect 295892 68546 295944 68552
rect 295996 19990 296024 70314
rect 295984 19984 296036 19990
rect 295984 19926 296036 19932
rect 296640 11898 296668 71726
rect 297284 69086 297312 71726
rect 297928 71726 297964 71754
rect 298634 71754 298662 72012
rect 299331 71754 299359 72012
rect 298634 71726 298692 71754
rect 297272 69080 297324 69086
rect 297272 69022 297324 69028
rect 296628 11892 296680 11898
rect 296628 11834 296680 11840
rect 294892 6886 295288 6914
rect 290188 6724 290240 6730
rect 290188 6666 290240 6672
rect 289084 6452 289136 6458
rect 289084 6394 289136 6400
rect 288992 6384 289044 6390
rect 288992 6326 289044 6332
rect 287796 3120 287848 3126
rect 287796 3062 287848 3068
rect 287808 480 287836 3062
rect 289004 480 289032 6326
rect 290200 480 290228 6666
rect 293684 6656 293736 6662
rect 293684 6598 293736 6604
rect 292580 6316 292632 6322
rect 292580 6258 292632 6264
rect 291384 2984 291436 2990
rect 291384 2926 291436 2932
rect 291396 480 291424 2926
rect 292592 480 292620 6258
rect 293696 480 293724 6598
rect 294892 480 294920 6886
rect 297272 6588 297324 6594
rect 297272 6530 297324 6536
rect 296076 6248 296128 6254
rect 296076 6190 296128 6196
rect 296088 480 296116 6190
rect 297284 480 297312 6530
rect 297928 5778 297956 71726
rect 298664 69086 298692 71726
rect 299216 71726 299359 71754
rect 300029 71754 300057 72012
rect 300727 71754 300755 72012
rect 301425 71754 301453 72012
rect 302123 71754 302151 72012
rect 302820 71754 302848 72012
rect 303518 71754 303546 72012
rect 300029 71726 300072 71754
rect 300727 71726 300808 71754
rect 298008 69080 298060 69086
rect 298008 69022 298060 69028
rect 298652 69080 298704 69086
rect 298652 69022 298704 69028
rect 297916 5772 297968 5778
rect 297916 5714 297968 5720
rect 298020 5710 298048 69022
rect 299216 5914 299244 71726
rect 299388 70372 299440 70378
rect 299388 70314 299440 70320
rect 299296 69080 299348 69086
rect 299296 69022 299348 69028
rect 299204 5908 299256 5914
rect 299204 5850 299256 5856
rect 299308 5846 299336 69022
rect 299296 5840 299348 5846
rect 299296 5782 299348 5788
rect 298008 5704 298060 5710
rect 298008 5646 298060 5652
rect 299400 2990 299428 70314
rect 300044 69086 300072 71726
rect 300032 69080 300084 69086
rect 300032 69022 300084 69028
rect 300676 69080 300728 69086
rect 300676 69022 300728 69028
rect 300688 16574 300716 69022
rect 300596 16546 300716 16574
rect 299664 6180 299716 6186
rect 299664 6122 299716 6128
rect 298468 2984 298520 2990
rect 298468 2926 298520 2932
rect 299388 2984 299440 2990
rect 299388 2926 299440 2932
rect 298480 480 298508 2926
rect 299676 480 299704 6122
rect 300596 5982 300624 16546
rect 300780 6914 300808 71726
rect 301424 71726 301453 71754
rect 302068 71726 302151 71754
rect 302804 71726 302848 71754
rect 303448 71726 303546 71754
rect 304216 71754 304244 72012
rect 304914 71754 304942 72012
rect 305612 71754 305640 72012
rect 306309 71754 306337 72012
rect 304216 71726 304304 71754
rect 304914 71726 304948 71754
rect 305612 71726 305684 71754
rect 301424 69086 301452 71726
rect 301412 69080 301464 69086
rect 301412 69022 301464 69028
rect 300688 6886 300808 6914
rect 300688 6050 300716 6886
rect 302068 6866 302096 71726
rect 302804 69086 302832 71726
rect 302148 69080 302200 69086
rect 302148 69022 302200 69028
rect 302792 69080 302844 69086
rect 302792 69022 302844 69028
rect 302056 6860 302108 6866
rect 302056 6802 302108 6808
rect 300768 6520 300820 6526
rect 300768 6462 300820 6468
rect 300676 6044 300728 6050
rect 300676 5986 300728 5992
rect 300584 5976 300636 5982
rect 300584 5918 300636 5924
rect 300780 480 300808 6462
rect 302160 6118 302188 69022
rect 303160 12300 303212 12306
rect 303160 12242 303212 12248
rect 302148 6112 302200 6118
rect 302148 6054 302200 6060
rect 301964 2984 302016 2990
rect 301964 2926 302016 2932
rect 301976 480 302004 2926
rect 303172 480 303200 12242
rect 303448 6730 303476 71726
rect 304276 69086 304304 71726
rect 303528 69080 303580 69086
rect 303528 69022 303580 69028
rect 304264 69080 304316 69086
rect 304264 69022 304316 69028
rect 304816 69080 304868 69086
rect 304816 69022 304868 69028
rect 303540 6798 303568 69022
rect 304356 9512 304408 9518
rect 304356 9454 304408 9460
rect 303528 6792 303580 6798
rect 303528 6734 303580 6740
rect 303436 6724 303488 6730
rect 303436 6666 303488 6672
rect 304368 480 304396 9454
rect 304828 6662 304856 69022
rect 304816 6656 304868 6662
rect 304816 6598 304868 6604
rect 304920 6594 304948 71726
rect 305656 69086 305684 71726
rect 306300 71726 306337 71754
rect 307007 71754 307035 72012
rect 307705 71754 307733 72012
rect 307007 71726 307064 71754
rect 305644 69080 305696 69086
rect 305644 69022 305696 69028
rect 306196 69080 306248 69086
rect 306196 69022 306248 69028
rect 304908 6588 304960 6594
rect 304908 6530 304960 6536
rect 306208 6526 306236 69022
rect 306196 6520 306248 6526
rect 306196 6462 306248 6468
rect 306300 6458 306328 71726
rect 307036 69086 307064 71726
rect 307588 71726 307733 71754
rect 308403 71754 308431 72012
rect 309101 71754 309129 72012
rect 309798 71754 309826 72012
rect 308403 71726 308444 71754
rect 307024 69080 307076 69086
rect 307024 69022 307076 69028
rect 306748 13524 306800 13530
rect 306748 13466 306800 13472
rect 306288 6452 306340 6458
rect 306288 6394 306340 6400
rect 305552 2916 305604 2922
rect 305552 2858 305604 2864
rect 305564 480 305592 2858
rect 306760 480 306788 13466
rect 307588 6322 307616 71726
rect 308416 69086 308444 71726
rect 308968 71726 309129 71754
rect 309796 71726 309826 71754
rect 310496 71754 310524 72012
rect 311194 71754 311222 72012
rect 310496 71726 310560 71754
rect 307668 69080 307720 69086
rect 307668 69022 307720 69028
rect 308404 69080 308456 69086
rect 308404 69022 308456 69028
rect 307680 6390 307708 69022
rect 308968 9654 308996 71726
rect 309796 69086 309824 71726
rect 310152 69624 310204 69630
rect 310152 69566 310204 69572
rect 309876 69284 309928 69290
rect 309876 69226 309928 69232
rect 309048 69080 309100 69086
rect 309048 69022 309100 69028
rect 309784 69080 309836 69086
rect 309784 69022 309836 69028
rect 308956 9648 309008 9654
rect 308956 9590 309008 9596
rect 307944 9308 307996 9314
rect 307944 9250 307996 9256
rect 307668 6384 307720 6390
rect 307668 6326 307720 6332
rect 307576 6316 307628 6322
rect 307576 6258 307628 6264
rect 307956 480 307984 9250
rect 309060 6254 309088 69022
rect 309888 64874 309916 69226
rect 310164 67182 310192 69566
rect 310336 69420 310388 69426
rect 310336 69362 310388 69368
rect 310348 68678 310376 69362
rect 310532 69154 310560 71726
rect 311176 71726 311222 71754
rect 311892 71754 311920 72012
rect 312590 71754 312618 72012
rect 311892 71726 311940 71754
rect 310520 69148 310572 69154
rect 310520 69090 310572 69096
rect 311176 69086 311204 71726
rect 311808 69148 311860 69154
rect 311808 69090 311860 69096
rect 310428 69080 310480 69086
rect 310428 69022 310480 69028
rect 311164 69080 311216 69086
rect 311164 69022 311216 69028
rect 311716 69080 311768 69086
rect 311716 69022 311768 69028
rect 310336 68672 310388 68678
rect 310336 68614 310388 68620
rect 310152 67176 310204 67182
rect 310152 67118 310204 67124
rect 309796 64846 309916 64874
rect 309796 15978 309824 64846
rect 309784 15972 309836 15978
rect 309784 15914 309836 15920
rect 310244 14748 310296 14754
rect 310244 14690 310296 14696
rect 309048 6248 309100 6254
rect 309048 6190 309100 6196
rect 309048 2848 309100 2854
rect 309048 2790 309100 2796
rect 309060 480 309088 2790
rect 310256 480 310284 14690
rect 310440 6186 310468 69022
rect 311728 9314 311756 69022
rect 311820 9518 311848 69090
rect 311912 69086 311940 71726
rect 312556 71726 312618 71754
rect 313287 71754 313315 72012
rect 313985 71754 314013 72012
rect 313287 71726 313320 71754
rect 311900 69080 311952 69086
rect 311900 69022 311952 69028
rect 312556 68338 312584 71726
rect 313188 69624 313240 69630
rect 313188 69566 313240 69572
rect 313096 69080 313148 69086
rect 313096 69022 313148 69028
rect 312544 68332 312596 68338
rect 312544 68274 312596 68280
rect 311808 9512 311860 9518
rect 311808 9454 311860 9460
rect 311716 9308 311768 9314
rect 311716 9250 311768 9256
rect 313108 9246 313136 69022
rect 311440 9240 311492 9246
rect 311440 9182 311492 9188
rect 313096 9240 313148 9246
rect 313096 9182 313148 9188
rect 310428 6180 310480 6186
rect 310428 6122 310480 6128
rect 311452 480 311480 9182
rect 313200 3602 313228 69566
rect 313292 18630 313320 71726
rect 313476 71726 314013 71754
rect 314683 71754 314711 72012
rect 315381 71754 315409 72012
rect 316079 71754 316107 72012
rect 316776 71754 316804 72012
rect 314683 71726 314884 71754
rect 313280 18624 313332 18630
rect 313280 18566 313332 18572
rect 313476 16114 313504 71726
rect 314752 68332 314804 68338
rect 314752 68274 314804 68280
rect 313464 16108 313516 16114
rect 313464 16050 313516 16056
rect 313832 12232 313884 12238
rect 313832 12174 313884 12180
rect 312636 3596 312688 3602
rect 312636 3538 312688 3544
rect 313188 3596 313240 3602
rect 313188 3538 313240 3544
rect 312648 480 312676 3538
rect 313844 480 313872 12174
rect 314764 3505 314792 68274
rect 314750 3496 314806 3505
rect 314750 3431 314806 3440
rect 314856 3369 314884 71726
rect 315316 71726 315409 71754
rect 316052 71726 316107 71754
rect 316420 71726 316804 71754
rect 317474 71754 317502 72012
rect 318172 71754 318200 72012
rect 317474 71726 317552 71754
rect 315316 68338 315344 71726
rect 315304 68332 315356 68338
rect 315304 68274 315356 68280
rect 315028 8424 315080 8430
rect 315028 8366 315080 8372
rect 314842 3360 314898 3369
rect 314842 3295 314898 3304
rect 315040 480 315068 8366
rect 316052 3466 316080 71726
rect 316316 16040 316368 16046
rect 316316 15982 316368 15988
rect 316132 3732 316184 3738
rect 316132 3674 316184 3680
rect 316144 3466 316172 3674
rect 316224 3596 316276 3602
rect 316224 3538 316276 3544
rect 316040 3460 316092 3466
rect 316040 3402 316092 3408
rect 316132 3460 316184 3466
rect 316132 3402 316184 3408
rect 316236 480 316264 3538
rect 316328 3482 316356 15982
rect 316420 3738 316448 71726
rect 316408 3732 316460 3738
rect 316408 3674 316460 3680
rect 317524 3670 317552 71726
rect 317616 71726 318200 71754
rect 318870 71754 318898 72012
rect 319568 71754 319596 72012
rect 318870 71726 318932 71754
rect 317512 3664 317564 3670
rect 317512 3606 317564 3612
rect 317616 3534 317644 71726
rect 318524 8492 318576 8498
rect 318524 8434 318576 8440
rect 317604 3528 317656 3534
rect 316328 3454 317368 3482
rect 317604 3470 317656 3476
rect 317340 480 317368 3454
rect 318536 480 318564 8434
rect 318904 3466 318932 71726
rect 319548 71726 319596 71754
rect 320265 71754 320293 72012
rect 320963 71754 320991 72012
rect 320265 71726 320312 71754
rect 319548 69290 319576 71726
rect 320284 69494 320312 71726
rect 320376 71726 320991 71754
rect 321560 71800 321612 71806
rect 321560 71742 321612 71748
rect 321661 71754 321689 72012
rect 322359 71806 322387 72012
rect 322347 71800 322399 71806
rect 320272 69488 320324 69494
rect 320272 69430 320324 69436
rect 319536 69284 319588 69290
rect 319536 69226 319588 69232
rect 320180 68808 320232 68814
rect 320180 68750 320232 68756
rect 320192 16574 320220 68750
rect 320376 17338 320404 71726
rect 320364 17332 320416 17338
rect 320364 17274 320416 17280
rect 320192 16546 320956 16574
rect 319720 3664 319772 3670
rect 319720 3606 319772 3612
rect 318892 3460 318944 3466
rect 318892 3402 318944 3408
rect 319732 480 319760 3606
rect 320928 480 320956 16546
rect 321572 14822 321600 71742
rect 321661 71726 321692 71754
rect 323057 71754 323085 72012
rect 323754 71754 323782 72012
rect 322347 71742 322399 71748
rect 321664 17270 321692 71726
rect 323044 71726 323085 71754
rect 323136 71726 323782 71754
rect 324320 71800 324372 71806
rect 324452 71754 324480 72012
rect 325150 71806 325178 72012
rect 324320 71742 324372 71748
rect 323044 69562 323072 71726
rect 323032 69556 323084 69562
rect 323032 69498 323084 69504
rect 321652 17264 321704 17270
rect 321652 17206 321704 17212
rect 323136 16182 323164 71726
rect 324228 69556 324280 69562
rect 324228 69498 324280 69504
rect 323124 16176 323176 16182
rect 323124 16118 323176 16124
rect 321560 14816 321612 14822
rect 321560 14758 321612 14764
rect 322112 8560 322164 8566
rect 322112 8502 322164 8508
rect 322124 480 322152 8502
rect 324240 3466 324268 69498
rect 324332 14890 324360 71742
rect 324424 71726 324480 71754
rect 325138 71800 325190 71806
rect 325848 71754 325876 72012
rect 326546 71754 326574 72012
rect 325138 71742 325190 71748
rect 325804 71726 325876 71754
rect 326540 71726 326574 71754
rect 327080 71800 327132 71806
rect 327243 71754 327271 72012
rect 327941 71806 327969 72012
rect 327080 71742 327132 71748
rect 324424 17406 324452 71726
rect 325804 70310 325832 71726
rect 325792 70304 325844 70310
rect 325792 70246 325844 70252
rect 326540 67250 326568 71726
rect 326528 67244 326580 67250
rect 326528 67186 326580 67192
rect 324412 17400 324464 17406
rect 324412 17342 324464 17348
rect 327092 16250 327120 71742
rect 327184 71726 327271 71754
rect 327929 71800 327981 71806
rect 327929 71742 327981 71748
rect 328460 71800 328512 71806
rect 328639 71754 328667 72012
rect 329337 71806 329365 72012
rect 328460 71742 328512 71748
rect 327184 18698 327212 71726
rect 327724 69148 327776 69154
rect 327724 69090 327776 69096
rect 327172 18692 327224 18698
rect 327172 18634 327224 18640
rect 327080 16244 327132 16250
rect 327080 16186 327132 16192
rect 324320 14884 324372 14890
rect 324320 14826 324372 14832
rect 327736 13598 327764 69090
rect 328472 17474 328500 71742
rect 328564 71726 328667 71754
rect 329325 71800 329377 71806
rect 329325 71742 329377 71748
rect 329840 71800 329892 71806
rect 330035 71754 330063 72012
rect 330732 71806 330760 72012
rect 329840 71742 329892 71748
rect 328564 44878 328592 71726
rect 328552 44872 328604 44878
rect 328552 44814 328604 44820
rect 329852 18766 329880 71742
rect 329944 71726 330063 71754
rect 330720 71800 330772 71806
rect 330720 71742 330772 71748
rect 331220 71800 331272 71806
rect 331430 71754 331458 72012
rect 332128 71806 332156 72012
rect 331220 71742 331272 71748
rect 329944 22778 329972 71726
rect 329932 22772 329984 22778
rect 329932 22714 329984 22720
rect 329840 18760 329892 18766
rect 329840 18702 329892 18708
rect 328460 17468 328512 17474
rect 328460 17410 328512 17416
rect 331232 14958 331260 71742
rect 331416 71726 331458 71754
rect 332116 71800 332168 71806
rect 332826 71754 332854 72012
rect 332116 71742 332168 71748
rect 332796 71726 332854 71754
rect 333524 71754 333552 72012
rect 333980 71800 334032 71806
rect 333524 71726 333560 71754
rect 334221 71754 334249 72012
rect 334919 71806 334947 72012
rect 333980 71742 334032 71748
rect 331312 47592 331364 47598
rect 331312 47534 331364 47540
rect 331324 16574 331352 47534
rect 331416 25566 331444 71726
rect 332796 69154 332824 71726
rect 332784 69148 332836 69154
rect 332784 69090 332836 69096
rect 333532 69086 333560 71726
rect 331864 69080 331916 69086
rect 331864 69022 331916 69028
rect 333520 69080 333572 69086
rect 333520 69022 333572 69028
rect 331876 50386 331904 69022
rect 331864 50380 331916 50386
rect 331864 50322 331916 50328
rect 331404 25560 331456 25566
rect 331404 25502 331456 25508
rect 331324 16546 331628 16574
rect 331220 14952 331272 14958
rect 331220 14894 331272 14900
rect 327724 13592 327776 13598
rect 327724 13534 327776 13540
rect 324412 13456 324464 13462
rect 324412 13398 324464 13404
rect 323308 3460 323360 3466
rect 323308 3402 323360 3408
rect 324228 3460 324280 3466
rect 324228 3402 324280 3408
rect 323320 480 323348 3402
rect 324424 480 324452 13398
rect 328000 13388 328052 13394
rect 328000 13330 328052 13336
rect 325608 8628 325660 8634
rect 325608 8570 325660 8576
rect 325620 480 325648 8570
rect 326804 3596 326856 3602
rect 326804 3538 326856 3544
rect 326816 480 326844 3538
rect 328012 480 328040 13330
rect 329196 8696 329248 8702
rect 329196 8638 329248 8644
rect 329208 480 329236 8638
rect 330392 3664 330444 3670
rect 330392 3606 330444 3612
rect 330404 480 330432 3606
rect 331600 480 331628 16546
rect 332692 8764 332744 8770
rect 332692 8706 332744 8712
rect 332704 480 332732 8706
rect 333888 3732 333940 3738
rect 333888 3674 333940 3680
rect 333900 480 333928 3674
rect 333992 3641 334020 71742
rect 334084 71726 334249 71754
rect 334907 71800 334959 71806
rect 334907 71742 334959 71748
rect 335452 71800 335504 71806
rect 335617 71754 335645 72012
rect 336315 71806 336343 72012
rect 335452 71742 335504 71748
rect 334084 17610 334112 71726
rect 334072 17604 334124 17610
rect 334072 17546 334124 17552
rect 335084 14680 335136 14686
rect 335084 14622 335136 14628
rect 333978 3632 334034 3641
rect 333978 3567 334034 3576
rect 335096 480 335124 14622
rect 335464 3806 335492 71742
rect 335556 71726 335645 71754
rect 336303 71800 336355 71806
rect 337013 71754 337041 72012
rect 337710 71754 337738 72012
rect 336303 71742 336355 71748
rect 336752 71726 337041 71754
rect 337120 71726 337738 71754
rect 338120 71800 338172 71806
rect 338120 71742 338172 71748
rect 335452 3800 335504 3806
rect 335556 3777 335584 71726
rect 336280 8832 336332 8838
rect 336280 8774 336332 8780
rect 335452 3742 335504 3748
rect 335542 3768 335598 3777
rect 335542 3703 335598 3712
rect 336292 480 336320 8774
rect 336752 3874 336780 71726
rect 337120 64874 337148 71726
rect 338028 70304 338080 70310
rect 338028 70246 338080 70252
rect 336844 64846 337148 64874
rect 336844 3942 336872 64846
rect 336832 3936 336884 3942
rect 336832 3878 336884 3884
rect 336740 3868 336792 3874
rect 336740 3810 336792 3816
rect 338040 3398 338068 70246
rect 338132 4078 338160 71742
rect 338304 49020 338356 49026
rect 338304 48962 338356 48968
rect 338120 4072 338172 4078
rect 338120 4014 338172 4020
rect 338316 3482 338344 48962
rect 338408 4010 338436 72012
rect 339106 71806 339134 72012
rect 339094 71800 339146 71806
rect 339804 71754 339832 72012
rect 340502 71754 340530 72012
rect 339094 71742 339146 71748
rect 339604 71726 339832 71754
rect 339880 71726 340530 71754
rect 340972 71800 341024 71806
rect 341199 71754 341227 72012
rect 341897 71806 341925 72012
rect 342595 71890 342623 72012
rect 342364 71862 342623 71890
rect 340972 71742 341024 71748
rect 339604 4146 339632 71726
rect 339880 64874 339908 71726
rect 339696 64846 339908 64874
rect 339592 4140 339644 4146
rect 339592 4082 339644 4088
rect 338396 4004 338448 4010
rect 338396 3946 338448 3952
rect 338316 3454 338712 3482
rect 337476 3392 337528 3398
rect 337476 3334 337528 3340
rect 338028 3392 338080 3398
rect 338028 3334 338080 3340
rect 337488 480 337516 3334
rect 338684 480 338712 3454
rect 339696 3330 339724 64846
rect 339868 8900 339920 8906
rect 339868 8842 339920 8848
rect 339684 3324 339736 3330
rect 339684 3266 339736 3272
rect 339880 480 339908 8842
rect 340984 6914 341012 71742
rect 341168 71726 341227 71754
rect 341885 71800 341937 71806
rect 341885 71742 341937 71748
rect 341064 11960 341116 11966
rect 341064 11902 341116 11908
rect 340892 6886 341012 6914
rect 340892 3262 340920 6886
rect 340972 3800 341024 3806
rect 340972 3742 341024 3748
rect 340880 3256 340932 3262
rect 340880 3198 340932 3204
rect 340984 480 341012 3742
rect 341076 3482 341104 11902
rect 341168 3874 341196 71726
rect 342364 70174 342392 71862
rect 343293 71754 343321 72012
rect 343991 71754 344019 72012
rect 344688 71754 344716 72012
rect 342456 71726 343321 71754
rect 343652 71726 344019 71754
rect 344204 71726 344716 71754
rect 345386 71754 345414 72012
rect 346084 71754 346112 72012
rect 346782 71754 346810 72012
rect 347480 71754 347508 72012
rect 348177 71754 348205 72012
rect 345386 71726 345428 71754
rect 342352 70168 342404 70174
rect 342352 70110 342404 70116
rect 342168 69488 342220 69494
rect 342168 69430 342220 69436
rect 342180 6914 342208 69430
rect 342352 19984 342404 19990
rect 342352 19926 342404 19932
rect 342088 6886 342208 6914
rect 341156 3868 341208 3874
rect 341156 3810 341208 3816
rect 342088 3806 342116 6886
rect 342076 3800 342128 3806
rect 342076 3742 342128 3748
rect 341076 3454 342208 3482
rect 342180 480 342208 3454
rect 342364 3074 342392 19926
rect 342456 3194 342484 71726
rect 342444 3188 342496 3194
rect 342444 3130 342496 3136
rect 343652 3126 343680 71726
rect 344204 64874 344232 71726
rect 345400 70242 345428 71726
rect 346044 71726 346112 71754
rect 346412 71726 346810 71754
rect 347424 71726 347508 71754
rect 347976 71726 348205 71754
rect 348875 71754 348903 72012
rect 349252 71800 349304 71806
rect 348875 71726 348924 71754
rect 349573 71754 349601 72012
rect 350271 71806 350299 72012
rect 350969 71890 350997 72012
rect 350644 71862 350997 71890
rect 349252 71742 349304 71748
rect 346044 70378 346072 71726
rect 346032 70372 346084 70378
rect 346032 70314 346084 70320
rect 345388 70236 345440 70242
rect 345388 70178 345440 70184
rect 345020 68740 345072 68746
rect 345020 68682 345072 68688
rect 343744 64846 344232 64874
rect 343640 3120 343692 3126
rect 342364 3046 343404 3074
rect 343640 3062 343692 3068
rect 343744 3058 343772 64846
rect 345032 16574 345060 68682
rect 345032 16546 345796 16574
rect 344560 4072 344612 4078
rect 344560 4014 344612 4020
rect 343376 480 343404 3046
rect 343732 3052 343784 3058
rect 343732 2994 343784 3000
rect 344572 480 344600 4014
rect 345768 480 345796 16546
rect 346412 2990 346440 71726
rect 347424 64874 347452 71726
rect 346504 64846 347452 64874
rect 346400 2984 346452 2990
rect 346400 2926 346452 2932
rect 346504 2922 346532 64846
rect 346952 12436 347004 12442
rect 346952 12378 347004 12384
rect 346492 2916 346544 2922
rect 346492 2858 346544 2864
rect 346964 480 346992 12378
rect 347976 2854 348004 71726
rect 348896 69630 348924 71726
rect 348884 69624 348936 69630
rect 348884 69566 348936 69572
rect 349264 16574 349292 71742
rect 349172 16546 349292 16574
rect 349448 71726 349601 71754
rect 350259 71800 350311 71806
rect 350259 71742 350311 71748
rect 348056 3596 348108 3602
rect 348056 3538 348108 3544
rect 347964 2848 348016 2854
rect 347964 2790 348016 2796
rect 348068 480 348096 3538
rect 349172 3534 349200 16546
rect 349344 15020 349396 15026
rect 349344 14962 349396 14968
rect 349252 13320 349304 13326
rect 349252 13262 349304 13268
rect 349160 3528 349212 3534
rect 349160 3470 349212 3476
rect 349264 480 349292 13262
rect 349356 3482 349384 14962
rect 349448 3942 349476 71726
rect 350644 69562 350672 71862
rect 351666 71754 351694 72012
rect 352364 71754 352392 72012
rect 353062 71754 353090 72012
rect 350736 71726 351694 71754
rect 351932 71726 352392 71754
rect 352484 71726 353090 71754
rect 353760 71754 353788 72012
rect 354458 71754 354486 72012
rect 355155 71754 355183 72012
rect 355853 71754 355881 72012
rect 356551 71754 356579 72012
rect 357249 71754 357277 72012
rect 357947 71754 357975 72012
rect 353760 71726 353800 71754
rect 350632 69556 350684 69562
rect 350632 69498 350684 69504
rect 349436 3936 349488 3942
rect 349436 3878 349488 3884
rect 350736 3670 350764 71726
rect 351932 3806 351960 71726
rect 352484 64874 352512 71726
rect 353772 70310 353800 71726
rect 354416 71726 354486 71754
rect 354692 71726 355183 71754
rect 355244 71726 355881 71754
rect 356164 71726 356579 71754
rect 356992 71726 357277 71754
rect 357452 71726 357975 71754
rect 358644 71754 358672 72012
rect 359342 71754 359370 72012
rect 360040 71754 360068 72012
rect 358644 71726 358768 71754
rect 359342 71726 359412 71754
rect 353760 70304 353812 70310
rect 353760 70246 353812 70252
rect 353944 69964 353996 69970
rect 353944 69906 353996 69912
rect 352024 64846 352512 64874
rect 352024 4010 352052 64846
rect 352840 14612 352892 14618
rect 352840 14554 352892 14560
rect 352012 4004 352064 4010
rect 352012 3946 352064 3952
rect 351920 3800 351972 3806
rect 351920 3742 351972 3748
rect 350724 3664 350776 3670
rect 350724 3606 350776 3612
rect 349356 3454 350488 3482
rect 350460 480 350488 3454
rect 351644 2984 351696 2990
rect 351644 2926 351696 2932
rect 351656 480 351684 2926
rect 352852 480 352880 14554
rect 353956 11966 353984 69906
rect 354416 69494 354444 71726
rect 354404 69488 354456 69494
rect 354404 69430 354456 69436
rect 354036 21412 354088 21418
rect 354036 21354 354088 21360
rect 353944 11960 353996 11966
rect 353944 11902 353996 11908
rect 354048 6914 354076 21354
rect 354128 16380 354180 16386
rect 354128 16322 354180 16328
rect 353956 6886 354076 6914
rect 353956 3670 353984 6886
rect 354036 4276 354088 4282
rect 354036 4218 354088 4224
rect 353944 3664 353996 3670
rect 353944 3606 353996 3612
rect 354048 480 354076 4218
rect 354140 3466 354168 16322
rect 354692 4078 354720 71726
rect 355244 64874 355272 71726
rect 354784 64846 355272 64874
rect 354680 4072 354732 4078
rect 354680 4014 354732 4020
rect 354784 3602 354812 64846
rect 354772 3596 354824 3602
rect 354772 3538 354824 3544
rect 355232 3528 355284 3534
rect 355232 3470 355284 3476
rect 354128 3460 354180 3466
rect 354128 3402 354180 3408
rect 355244 480 355272 3470
rect 356164 2990 356192 71726
rect 356992 64874 357020 71726
rect 356256 64846 357020 64874
rect 356256 3534 356284 64846
rect 356336 7064 356388 7070
rect 356336 7006 356388 7012
rect 356244 3528 356296 3534
rect 356244 3470 356296 3476
rect 356152 2984 356204 2990
rect 356152 2926 356204 2932
rect 356348 480 356376 7006
rect 357452 3534 357480 71726
rect 358740 6914 358768 71726
rect 359384 69086 359412 71726
rect 360028 71726 360068 71754
rect 360738 71754 360766 72012
rect 361436 71754 361464 72012
rect 362133 71754 362161 72012
rect 362831 71754 362859 72012
rect 363529 71754 363557 72012
rect 364227 71754 364255 72012
rect 364925 71754 364953 72012
rect 365622 71754 365650 72012
rect 360738 71726 360792 71754
rect 361436 71726 361528 71754
rect 362133 71726 362172 71754
rect 359372 69080 359424 69086
rect 359372 69022 359424 69028
rect 359924 7132 359976 7138
rect 359924 7074 359976 7080
rect 358648 6886 358768 6914
rect 357532 3664 357584 3670
rect 357532 3606 357584 3612
rect 357440 3528 357492 3534
rect 357440 3470 357492 3476
rect 357544 480 357572 3606
rect 358648 3602 358676 6886
rect 358636 3596 358688 3602
rect 358636 3538 358688 3544
rect 358728 3528 358780 3534
rect 358728 3470 358780 3476
rect 358740 480 358768 3470
rect 359936 480 359964 7074
rect 360028 3670 360056 71726
rect 360764 69086 360792 71726
rect 360108 69080 360160 69086
rect 360108 69022 360160 69028
rect 360752 69080 360804 69086
rect 360752 69022 360804 69028
rect 361396 69080 361448 69086
rect 361396 69022 361448 69028
rect 360016 3664 360068 3670
rect 360016 3606 360068 3612
rect 360120 3194 360148 69022
rect 360844 13728 360896 13734
rect 360844 13670 360896 13676
rect 360856 3942 360884 13670
rect 361408 4146 361436 69022
rect 361396 4140 361448 4146
rect 361396 4082 361448 4088
rect 361500 4010 361528 71726
rect 362144 69086 362172 71726
rect 362788 71726 362859 71754
rect 363524 71726 363557 71754
rect 364168 71726 364255 71754
rect 364904 71726 364953 71754
rect 365548 71726 365650 71754
rect 366320 71754 366348 72012
rect 367018 71754 367046 72012
rect 367716 71754 367744 72012
rect 368414 71754 368442 72012
rect 366320 71726 366404 71754
rect 367018 71726 367048 71754
rect 367716 71726 367784 71754
rect 362132 69080 362184 69086
rect 362132 69022 362184 69028
rect 361488 4004 361540 4010
rect 361488 3946 361540 3952
rect 360844 3936 360896 3942
rect 360844 3878 360896 3884
rect 362788 3806 362816 71726
rect 363524 69086 363552 71726
rect 362868 69080 362920 69086
rect 362868 69022 362920 69028
rect 363512 69080 363564 69086
rect 363512 69022 363564 69028
rect 362880 3874 362908 69022
rect 363512 7200 363564 7206
rect 363512 7142 363564 7148
rect 362868 3868 362920 3874
rect 362868 3810 362920 3816
rect 362776 3800 362828 3806
rect 362776 3742 362828 3748
rect 362316 3596 362368 3602
rect 362316 3538 362368 3544
rect 361120 3460 361172 3466
rect 361120 3402 361172 3408
rect 360108 3188 360160 3194
rect 360108 3130 360160 3136
rect 361132 480 361160 3402
rect 362328 480 362356 3538
rect 363524 480 363552 7142
rect 364168 3670 364196 71726
rect 364904 69086 364932 71726
rect 364248 69080 364300 69086
rect 364248 69022 364300 69028
rect 364892 69080 364944 69086
rect 364892 69022 364944 69028
rect 364260 3738 364288 69022
rect 364616 3936 364668 3942
rect 364616 3878 364668 3884
rect 364248 3732 364300 3738
rect 364248 3674 364300 3680
rect 364156 3664 364208 3670
rect 364156 3606 364208 3612
rect 364628 480 364656 3878
rect 365548 3466 365576 71726
rect 366376 69086 366404 71726
rect 365628 69080 365680 69086
rect 365628 69022 365680 69028
rect 366364 69080 366416 69086
rect 366364 69022 366416 69028
rect 366916 69080 366968 69086
rect 366916 69022 366968 69028
rect 365640 3534 365668 69022
rect 366928 16574 366956 69022
rect 366836 16546 366956 16574
rect 365628 3528 365680 3534
rect 365628 3470 365680 3476
rect 365536 3460 365588 3466
rect 365536 3402 365588 3408
rect 366836 3330 366864 16546
rect 367020 11778 367048 71726
rect 367756 69358 367784 71726
rect 368400 71726 368442 71754
rect 369111 71754 369139 72012
rect 369809 71754 369837 72012
rect 369111 71726 369164 71754
rect 367744 69352 367796 69358
rect 367744 69294 367796 69300
rect 367100 17536 367152 17542
rect 367100 17478 367152 17484
rect 367112 16574 367140 17478
rect 367112 16546 368244 16574
rect 366928 11750 367048 11778
rect 366824 3324 366876 3330
rect 366824 3266 366876 3272
rect 365812 3188 365864 3194
rect 365812 3130 365864 3136
rect 365824 480 365852 3130
rect 366928 2854 366956 11750
rect 367008 7268 367060 7274
rect 367008 7210 367060 7216
rect 366916 2848 366968 2854
rect 366916 2790 366968 2796
rect 367020 480 367048 7210
rect 368216 480 368244 16546
rect 368400 2922 368428 71726
rect 369136 69086 369164 71726
rect 369780 71726 369837 71754
rect 370507 71754 370535 72012
rect 371205 71754 371233 72012
rect 371903 71754 371931 72012
rect 370507 71726 370544 71754
rect 369124 69080 369176 69086
rect 369124 69022 369176 69028
rect 369676 69080 369728 69086
rect 369676 69022 369728 69028
rect 369400 3596 369452 3602
rect 369400 3538 369452 3544
rect 368388 2916 368440 2922
rect 368388 2858 368440 2864
rect 369412 480 369440 3538
rect 369688 2990 369716 69022
rect 369780 3058 369808 71726
rect 370516 69426 370544 71726
rect 371160 71726 371233 71754
rect 371896 71726 371931 71754
rect 372600 71754 372628 72012
rect 373298 71754 373326 72012
rect 372600 71726 372660 71754
rect 370504 69420 370556 69426
rect 370504 69362 370556 69368
rect 370596 7336 370648 7342
rect 370596 7278 370648 7284
rect 369768 3052 369820 3058
rect 369768 2994 369820 3000
rect 369676 2984 369728 2990
rect 369676 2926 369728 2932
rect 370608 480 370636 7278
rect 371160 3126 371188 71726
rect 371792 69692 371844 69698
rect 371792 69634 371844 69640
rect 371804 64874 371832 69634
rect 371896 69494 371924 71726
rect 372632 69562 372660 71726
rect 373276 71726 373326 71754
rect 373996 71754 374024 72012
rect 374694 71754 374722 72012
rect 373996 71726 374040 71754
rect 374694 71726 374776 71754
rect 372620 69556 372672 69562
rect 372620 69498 372672 69504
rect 371884 69488 371936 69494
rect 371884 69430 371936 69436
rect 373276 69086 373304 71726
rect 374012 69630 374040 71726
rect 374000 69624 374052 69630
rect 374000 69566 374052 69572
rect 374748 69086 374776 71726
rect 375392 70378 375420 72012
rect 376089 71754 376117 72012
rect 376787 71754 376815 72012
rect 376089 71726 376156 71754
rect 375380 70372 375432 70378
rect 375380 70314 375432 70320
rect 376128 69086 376156 71726
rect 376772 71726 376815 71754
rect 377485 71754 377513 72012
rect 378183 71754 378211 72012
rect 378881 71754 378909 72012
rect 379578 71754 379606 72012
rect 380276 71754 380304 72012
rect 377485 71726 377536 71754
rect 378183 71726 378272 71754
rect 378881 71726 378916 71754
rect 379578 71726 379652 71754
rect 376772 69698 376800 71726
rect 376760 69692 376812 69698
rect 376760 69634 376812 69640
rect 377508 69086 377536 71726
rect 378244 70310 378272 71726
rect 378232 70304 378284 70310
rect 378232 70246 378284 70252
rect 378888 69086 378916 71726
rect 379624 70174 379652 71726
rect 380268 71726 380304 71754
rect 380974 71754 381002 72012
rect 381672 71754 381700 72012
rect 380974 71726 381032 71754
rect 379612 70168 379664 70174
rect 379612 70110 379664 70116
rect 380268 69086 380296 71726
rect 381004 70242 381032 71726
rect 381648 71726 381700 71754
rect 382370 71754 382398 72012
rect 383067 71754 383095 72012
rect 383765 71754 383793 72012
rect 382370 71726 382412 71754
rect 383067 71726 383516 71754
rect 380992 70236 381044 70242
rect 380992 70178 381044 70184
rect 381648 69086 381676 71726
rect 382384 69086 382412 71726
rect 373264 69080 373316 69086
rect 373264 69022 373316 69028
rect 373908 69080 373960 69086
rect 373908 69022 373960 69028
rect 374736 69080 374788 69086
rect 374736 69022 374788 69028
rect 375288 69080 375340 69086
rect 375288 69022 375340 69028
rect 376116 69080 376168 69086
rect 376116 69022 376168 69028
rect 376668 69080 376720 69086
rect 376668 69022 376720 69028
rect 377496 69080 377548 69086
rect 377496 69022 377548 69028
rect 378048 69080 378100 69086
rect 378048 69022 378100 69028
rect 378876 69080 378928 69086
rect 378876 69022 378928 69028
rect 379428 69080 379480 69086
rect 379428 69022 379480 69028
rect 380256 69080 380308 69086
rect 380256 69022 380308 69028
rect 380808 69080 380860 69086
rect 380808 69022 380860 69028
rect 381636 69080 381688 69086
rect 381636 69022 381688 69028
rect 382188 69080 382240 69086
rect 382188 69022 382240 69028
rect 382372 69080 382424 69086
rect 382372 69022 382424 69028
rect 371804 64846 371924 64874
rect 371700 16312 371752 16318
rect 371700 16254 371752 16260
rect 371148 3120 371200 3126
rect 371148 3062 371200 3068
rect 371712 480 371740 16254
rect 371896 7342 371924 64846
rect 371884 7336 371936 7342
rect 371884 7278 371936 7284
rect 372896 4140 372948 4146
rect 372896 4082 372948 4088
rect 372908 480 372936 4082
rect 373920 3194 373948 69022
rect 374000 67312 374052 67318
rect 374000 67254 374052 67260
rect 374012 3262 374040 67254
rect 374092 7404 374144 7410
rect 374092 7346 374144 7352
rect 374000 3256 374052 3262
rect 374000 3198 374052 3204
rect 373908 3188 373960 3194
rect 373908 3130 373960 3136
rect 374104 480 374132 7346
rect 375300 6914 375328 69022
rect 375208 6886 375328 6914
rect 375208 3330 375236 6886
rect 376484 4004 376536 4010
rect 376484 3946 376536 3952
rect 375196 3324 375248 3330
rect 375196 3266 375248 3272
rect 375288 3256 375340 3262
rect 375288 3198 375340 3204
rect 375300 480 375328 3198
rect 376496 480 376524 3946
rect 376680 3330 376708 69022
rect 377680 7472 377732 7478
rect 377680 7414 377732 7420
rect 376668 3324 376720 3330
rect 376668 3266 376720 3272
rect 377692 480 377720 7414
rect 378060 3398 378088 69022
rect 378876 9784 378928 9790
rect 378876 9726 378928 9732
rect 378048 3392 378100 3398
rect 378048 3334 378100 3340
rect 378888 480 378916 9726
rect 379440 4146 379468 69022
rect 379428 4140 379480 4146
rect 379428 4082 379480 4088
rect 380820 4078 380848 69022
rect 381176 7540 381228 7546
rect 381176 7482 381228 7488
rect 380808 4072 380860 4078
rect 380808 4014 380860 4020
rect 379980 3868 380032 3874
rect 379980 3810 380032 3816
rect 379992 480 380020 3810
rect 381188 480 381216 7482
rect 382200 4010 382228 69022
rect 383488 64394 383516 71726
rect 383764 71726 383793 71754
rect 384463 71754 384491 72012
rect 385161 71754 385189 72012
rect 384463 71726 384528 71754
rect 383764 69290 383792 71726
rect 383752 69284 383804 69290
rect 383752 69226 383804 69232
rect 383568 69080 383620 69086
rect 383568 69022 383620 69028
rect 383476 64388 383528 64394
rect 383476 64330 383528 64336
rect 383580 17270 383608 69022
rect 384500 68882 384528 71726
rect 385144 71726 385189 71754
rect 385859 71754 385887 72012
rect 386556 71754 386584 72012
rect 387254 71754 387282 72012
rect 387952 71754 387980 72012
rect 388650 71754 388678 72012
rect 385859 71726 385908 71754
rect 386556 71726 386644 71754
rect 387254 71726 387288 71754
rect 387952 71726 388024 71754
rect 384488 68876 384540 68882
rect 384488 68818 384540 68824
rect 385144 67318 385172 71726
rect 385880 69086 385908 71726
rect 385868 69080 385920 69086
rect 385868 69022 385920 69028
rect 386328 69080 386380 69086
rect 386328 69022 386380 69028
rect 385132 67312 385184 67318
rect 385132 67254 385184 67260
rect 386340 18630 386368 69022
rect 386616 68814 386644 71726
rect 386604 68808 386656 68814
rect 386604 68750 386656 68756
rect 387260 67250 387288 71726
rect 387248 67244 387300 67250
rect 387248 67186 387300 67192
rect 387996 65890 388024 71726
rect 388640 71726 388678 71754
rect 389348 71754 389376 72012
rect 390045 71754 390073 72012
rect 389348 71726 389404 71754
rect 388640 69086 388668 71726
rect 389376 69154 389404 71726
rect 390020 71726 390073 71754
rect 390743 71754 390771 72012
rect 391441 71754 391469 72012
rect 392139 71754 392167 72012
rect 390743 71726 390784 71754
rect 391441 71726 391520 71754
rect 389364 69148 389416 69154
rect 389364 69090 389416 69096
rect 390020 69086 390048 71726
rect 390756 69154 390784 71726
rect 390376 69148 390428 69154
rect 390376 69090 390428 69096
rect 390744 69148 390796 69154
rect 390744 69090 390796 69096
rect 388628 69080 388680 69086
rect 388628 69022 388680 69028
rect 389088 69080 389140 69086
rect 389088 69022 389140 69028
rect 390008 69080 390060 69086
rect 390008 69022 390060 69028
rect 387984 65884 388036 65890
rect 387984 65826 388036 65832
rect 389100 58682 389128 69022
rect 390388 64326 390416 69090
rect 390468 69080 390520 69086
rect 390468 69022 390520 69028
rect 390376 64320 390428 64326
rect 390376 64262 390428 64268
rect 389088 58676 389140 58682
rect 389088 58618 389140 58624
rect 390480 21418 390508 69022
rect 391492 68746 391520 71726
rect 392136 71726 392167 71754
rect 392837 71754 392865 72012
rect 393534 71754 393562 72012
rect 392837 71726 393268 71754
rect 392136 69086 392164 71726
rect 392400 69148 392452 69154
rect 392400 69090 392452 69096
rect 392124 69080 392176 69086
rect 392124 69022 392176 69028
rect 391480 68740 391532 68746
rect 391480 68682 391532 68688
rect 392412 65822 392440 69090
rect 393136 69080 393188 69086
rect 393136 69022 393188 69028
rect 392400 65816 392452 65822
rect 392400 65758 392452 65764
rect 393148 62898 393176 69022
rect 393136 62892 393188 62898
rect 393136 62834 393188 62840
rect 393240 22778 393268 71726
rect 393516 71726 393562 71754
rect 394232 71754 394260 72012
rect 394930 71754 394958 72012
rect 395628 71754 395656 72012
rect 396326 71754 396354 72012
rect 397023 71754 397051 72012
rect 397721 71754 397749 72012
rect 398419 71754 398447 72012
rect 399117 71754 399145 72012
rect 399815 71754 399843 72012
rect 400512 71754 400540 72012
rect 394232 71726 394648 71754
rect 394930 71726 395016 71754
rect 395628 71726 396028 71754
rect 396326 71726 396396 71754
rect 397023 71726 397408 71754
rect 397721 71726 397776 71754
rect 398419 71726 398696 71754
rect 399117 71726 399156 71754
rect 399815 71726 400076 71754
rect 393516 69086 393544 71726
rect 393504 69080 393556 69086
rect 393504 69022 393556 69028
rect 394516 69080 394568 69086
rect 394516 69022 394568 69028
rect 394528 64258 394556 69022
rect 394516 64252 394568 64258
rect 394516 64194 394568 64200
rect 394620 50386 394648 71726
rect 394988 69086 395016 71726
rect 394976 69080 395028 69086
rect 394976 69022 395028 69028
rect 395896 69080 395948 69086
rect 395896 69022 395948 69028
rect 395908 62830 395936 69022
rect 395896 62824 395948 62830
rect 395896 62766 395948 62772
rect 394608 50380 394660 50386
rect 394608 50322 394660 50328
rect 393228 22772 393280 22778
rect 393228 22714 393280 22720
rect 390468 21412 390520 21418
rect 390468 21354 390520 21360
rect 386328 18624 386380 18630
rect 386328 18566 386380 18572
rect 383568 17264 383620 17270
rect 383568 17206 383620 17212
rect 393044 10056 393096 10062
rect 393044 9998 393096 10004
rect 389456 9988 389508 9994
rect 389456 9930 389508 9936
rect 385960 9920 386012 9926
rect 385960 9862 386012 9868
rect 382372 9852 382424 9858
rect 382372 9794 382424 9800
rect 382188 4004 382240 4010
rect 382188 3946 382240 3952
rect 382384 480 382412 9794
rect 384764 8288 384816 8294
rect 384764 8230 384816 8236
rect 383568 3800 383620 3806
rect 383568 3742 383620 3748
rect 383580 480 383608 3742
rect 384776 480 384804 8230
rect 385972 480 386000 9862
rect 388260 8220 388312 8226
rect 388260 8162 388312 8168
rect 387156 3732 387208 3738
rect 387156 3674 387208 3680
rect 387168 480 387196 3674
rect 388272 480 388300 8162
rect 389468 480 389496 9930
rect 391848 8152 391900 8158
rect 391848 8094 391900 8100
rect 390652 3664 390704 3670
rect 390652 3606 390704 3612
rect 390664 480 390692 3606
rect 391860 480 391888 8094
rect 393056 480 393084 9998
rect 395344 8084 395396 8090
rect 395344 8026 395396 8032
rect 394240 3596 394292 3602
rect 394240 3538 394292 3544
rect 394252 480 394280 3538
rect 395356 480 395384 8026
rect 396000 3806 396028 71726
rect 396368 69086 396396 71726
rect 396356 69080 396408 69086
rect 396356 69022 396408 69028
rect 397276 69080 397328 69086
rect 397276 69022 397328 69028
rect 396540 10124 396592 10130
rect 396540 10066 396592 10072
rect 395988 3800 396040 3806
rect 395988 3742 396040 3748
rect 396552 480 396580 10066
rect 397288 3874 397316 69022
rect 397380 3942 397408 71726
rect 397748 69086 397776 71726
rect 397736 69080 397788 69086
rect 397736 69022 397788 69028
rect 397368 3936 397420 3942
rect 397368 3878 397420 3884
rect 397276 3868 397328 3874
rect 397276 3810 397328 3816
rect 398668 3670 398696 71726
rect 399128 69086 399156 71726
rect 398748 69080 398800 69086
rect 398748 69022 398800 69028
rect 399116 69080 399168 69086
rect 399116 69022 399168 69028
rect 398760 3738 398788 69022
rect 400048 16574 400076 71726
rect 400508 71726 400540 71754
rect 401210 71754 401238 72012
rect 401908 71754 401936 72012
rect 401210 71726 401456 71754
rect 400508 69086 400536 71726
rect 400128 69080 400180 69086
rect 400128 69022 400180 69028
rect 400496 69080 400548 69086
rect 400496 69022 400548 69028
rect 399956 16546 400076 16574
rect 398840 10192 398892 10198
rect 398840 10134 398892 10140
rect 398748 3732 398800 3738
rect 398748 3674 398800 3680
rect 398656 3664 398708 3670
rect 398656 3606 398708 3612
rect 398852 3534 398880 10134
rect 398932 8016 398984 8022
rect 398932 7958 398984 7964
rect 397736 3528 397788 3534
rect 397736 3470 397788 3476
rect 398840 3528 398892 3534
rect 398840 3470 398892 3476
rect 397748 480 397776 3470
rect 398944 480 398972 7958
rect 399956 3806 399984 16546
rect 400140 6914 400168 69022
rect 400048 6886 400168 6914
rect 399944 3800 399996 3806
rect 399944 3742 399996 3748
rect 400048 3602 400076 6886
rect 401428 3641 401456 71726
rect 401888 71726 401936 71754
rect 402606 71754 402634 72012
rect 402916 71754 402944 72012
rect 402606 71726 402836 71754
rect 401888 69086 401916 71726
rect 401508 69080 401560 69086
rect 401508 69022 401560 69028
rect 401876 69080 401928 69086
rect 401876 69022 401928 69028
rect 401414 3632 401470 3641
rect 400036 3596 400088 3602
rect 401414 3567 401470 3576
rect 400036 3538 400088 3544
rect 400128 3528 400180 3534
rect 400128 3470 400180 3476
rect 400140 480 400168 3470
rect 401520 3466 401548 69022
rect 402520 7948 402572 7954
rect 402520 7890 402572 7896
rect 401324 3460 401376 3466
rect 401324 3402 401376 3408
rect 401508 3460 401560 3466
rect 401508 3402 401560 3408
rect 401336 480 401364 3402
rect 402532 480 402560 7890
rect 402808 3505 402836 71726
rect 402900 71726 402944 71754
rect 403304 71754 403332 72012
rect 403304 71726 403388 71754
rect 402794 3496 402850 3505
rect 402794 3431 402850 3440
rect 402900 3369 402928 71726
rect 403360 69154 403388 71726
rect 403348 69148 403400 69154
rect 403348 69090 403400 69096
rect 404176 69148 404228 69154
rect 404176 69090 404228 69096
rect 404188 64874 404216 69090
rect 404268 69080 404320 69086
rect 404268 69022 404320 69028
rect 404280 68338 404308 69022
rect 404268 68332 404320 68338
rect 404268 68274 404320 68280
rect 404188 64846 404308 64874
rect 403624 10260 403676 10266
rect 403624 10202 403676 10208
rect 402886 3360 402942 3369
rect 402886 3295 402942 3304
rect 403636 480 403664 10202
rect 404280 3777 404308 64846
rect 406016 7880 406068 7886
rect 406016 7822 406068 7828
rect 404266 3768 404322 3777
rect 404266 3703 404322 3712
rect 404820 2848 404872 2854
rect 404820 2790 404872 2796
rect 404832 480 404860 2790
rect 406028 480 406056 7822
rect 406396 5642 406424 72791
rect 406488 20670 406516 77551
rect 406580 33114 406608 83263
rect 406672 46918 406700 88839
rect 406764 60722 406792 94551
rect 406856 73166 406884 100263
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 406844 73160 406896 73166
rect 406844 73102 406896 73108
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 447140 70372 447192 70378
rect 447140 70314 447192 70320
rect 410524 70100 410576 70106
rect 410524 70042 410576 70048
rect 407120 69352 407172 69358
rect 407120 69294 407172 69300
rect 406752 60716 406804 60722
rect 406752 60658 406804 60664
rect 406660 46912 406712 46918
rect 406660 46854 406712 46860
rect 406568 33108 406620 33114
rect 406568 33050 406620 33056
rect 406476 20664 406528 20670
rect 406476 20606 406528 20612
rect 406384 5636 406436 5642
rect 406384 5578 406436 5584
rect 407132 2922 407160 69294
rect 407212 11008 407264 11014
rect 407212 10950 407264 10956
rect 407120 2916 407172 2922
rect 407120 2858 407172 2864
rect 407224 480 407252 10950
rect 410536 7818 410564 70042
rect 418804 70032 418856 70038
rect 418804 69974 418856 69980
rect 413284 69828 413336 69834
rect 413284 69770 413336 69776
rect 411904 69760 411956 69766
rect 411904 69702 411956 69708
rect 410800 10940 410852 10946
rect 410800 10882 410852 10888
rect 409604 7812 409656 7818
rect 409604 7754 409656 7760
rect 410524 7812 410576 7818
rect 410524 7754 410576 7760
rect 408408 2916 408460 2922
rect 408408 2858 408460 2864
rect 408420 480 408448 2858
rect 409616 480 409644 7754
rect 410812 480 410840 10882
rect 411916 7886 411944 69702
rect 411904 7880 411956 7886
rect 411904 7822 411956 7828
rect 413296 7750 413324 69770
rect 414664 69284 414716 69290
rect 414664 69226 414716 69232
rect 414676 10878 414704 69226
rect 414296 10872 414348 10878
rect 414296 10814 414348 10820
rect 414664 10872 414716 10878
rect 414664 10814 414716 10820
rect 413100 7744 413152 7750
rect 413100 7686 413152 7692
rect 413284 7744 413336 7750
rect 413284 7686 413336 7692
rect 411904 2848 411956 2854
rect 411904 2790 411956 2796
rect 411916 480 411944 2790
rect 413112 480 413140 7686
rect 414308 480 414336 10814
rect 417884 10804 417936 10810
rect 417884 10746 417936 10752
rect 416688 7676 416740 7682
rect 416688 7618 416740 7624
rect 415492 2984 415544 2990
rect 415492 2926 415544 2932
rect 415504 480 415532 2926
rect 416700 480 416728 7618
rect 417896 480 417924 10746
rect 418816 7682 418844 69974
rect 440240 69624 440292 69630
rect 440240 69566 440292 69572
rect 431960 69556 432012 69562
rect 431960 69498 432012 69504
rect 429200 69488 429252 69494
rect 429200 69430 429252 69436
rect 422300 69420 422352 69426
rect 422300 69362 422352 69368
rect 422312 16574 422340 69362
rect 423680 67040 423732 67046
rect 423680 66982 423732 66988
rect 423692 16574 423720 66982
rect 429212 16574 429240 69430
rect 430580 68536 430632 68542
rect 430580 68478 430632 68484
rect 430592 16574 430620 68478
rect 422312 16546 422616 16574
rect 423692 16546 423812 16574
rect 429212 16546 429700 16574
rect 430592 16546 430896 16574
rect 421380 10736 421432 10742
rect 421380 10678 421432 10684
rect 418804 7676 418856 7682
rect 418804 7618 418856 7624
rect 420184 7608 420236 7614
rect 420184 7550 420236 7556
rect 418988 3052 419040 3058
rect 418988 2994 419040 3000
rect 419000 480 419028 2994
rect 420196 480 420224 7550
rect 421392 480 421420 10678
rect 422588 480 422616 16546
rect 423784 480 423812 16546
rect 427268 11960 427320 11966
rect 427268 11902 427320 11908
rect 424968 10668 425020 10674
rect 424968 10610 425020 10616
rect 424980 480 425008 10610
rect 426164 3120 426216 3126
rect 426164 3062 426216 3068
rect 426176 480 426204 3062
rect 427280 480 427308 11902
rect 428464 10600 428516 10606
rect 428464 10542 428516 10548
rect 428476 480 428504 10542
rect 429672 480 429700 16546
rect 430868 480 430896 16546
rect 431972 3126 432000 69498
rect 440252 16574 440280 69566
rect 447152 16574 447180 70314
rect 454040 70304 454092 70310
rect 454040 70246 454092 70252
rect 448520 65612 448572 65618
rect 448520 65554 448572 65560
rect 448532 16574 448560 65554
rect 454052 16574 454080 70246
rect 460940 70236 460992 70242
rect 460940 70178 460992 70184
rect 456892 64184 456944 64190
rect 456892 64126 456944 64132
rect 440252 16546 440372 16574
rect 447152 16546 447456 16574
rect 448532 16546 448652 16574
rect 454052 16546 454540 16574
rect 437940 14476 437992 14482
rect 437940 14418 437992 14424
rect 434444 13252 434496 13258
rect 434444 13194 434496 13200
rect 432052 10532 432104 10538
rect 432052 10474 432104 10480
rect 431960 3120 432012 3126
rect 431960 3062 432012 3068
rect 432064 480 432092 10474
rect 433248 3120 433300 3126
rect 433248 3062 433300 3068
rect 433260 480 433288 3062
rect 434456 480 434484 13194
rect 435548 10464 435600 10470
rect 435548 10406 435600 10412
rect 435560 480 435588 10406
rect 436744 3188 436796 3194
rect 436744 3130 436796 3136
rect 436756 480 436784 3130
rect 437952 480 437980 14418
rect 439136 10396 439188 10402
rect 439136 10338 439188 10344
rect 439148 480 439176 10338
rect 440344 480 440372 16546
rect 441528 15904 441580 15910
rect 441528 15846 441580 15852
rect 441540 480 441568 15846
rect 446220 12164 446272 12170
rect 446220 12106 446272 12112
rect 445024 11824 445076 11830
rect 445024 11766 445076 11772
rect 442632 10328 442684 10334
rect 442632 10270 442684 10276
rect 442644 480 442672 10270
rect 443828 3256 443880 3262
rect 443828 3198 443880 3204
rect 443840 480 443868 3198
rect 445036 480 445064 11766
rect 446232 480 446260 12106
rect 447428 480 447456 16546
rect 448624 480 448652 16546
rect 452108 13184 452160 13190
rect 452108 13126 452160 13132
rect 449808 12096 449860 12102
rect 449808 12038 449860 12044
rect 449820 480 449848 12038
rect 450912 3324 450964 3330
rect 450912 3266 450964 3272
rect 450924 480 450952 3266
rect 452120 480 452148 13126
rect 453304 12028 453356 12034
rect 453304 11970 453356 11976
rect 453316 480 453344 11970
rect 454512 480 454540 16546
rect 455696 9580 455748 9586
rect 455696 9522 455748 9528
rect 455708 480 455736 9522
rect 456904 480 456932 64126
rect 459560 24132 459612 24138
rect 459560 24074 459612 24080
rect 459572 16574 459600 24074
rect 460952 16574 460980 70178
rect 467840 70168 467892 70174
rect 467840 70110 467892 70116
rect 466460 67108 466512 67114
rect 466460 67050 466512 67056
rect 463700 65748 463752 65754
rect 463700 65690 463752 65696
rect 463712 16574 463740 65690
rect 466472 16574 466500 67050
rect 467852 16574 467880 70110
rect 474740 69964 474792 69970
rect 474740 69906 474792 69912
rect 472624 69896 472676 69902
rect 472624 69838 472676 69844
rect 470600 65680 470652 65686
rect 470600 65622 470652 65628
rect 470612 16574 470640 65622
rect 459572 16546 460428 16574
rect 460952 16546 461624 16574
rect 463712 16546 464016 16574
rect 466472 16546 467512 16574
rect 467852 16546 468708 16574
rect 470612 16546 471100 16574
rect 459192 9444 459244 9450
rect 459192 9386 459244 9392
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 9386
rect 460400 480 460428 16546
rect 461596 480 461624 16546
rect 462780 9376 462832 9382
rect 462780 9318 462832 9324
rect 462792 480 462820 9318
rect 463988 480 464016 16546
rect 466276 9172 466328 9178
rect 466276 9114 466328 9120
rect 465172 4140 465224 4146
rect 465172 4082 465224 4088
rect 465184 480 465212 4082
rect 466288 480 466316 9114
rect 467484 480 467512 16546
rect 468680 480 468708 16546
rect 469864 9104 469916 9110
rect 469864 9046 469916 9052
rect 469876 480 469904 9046
rect 471072 480 471100 16546
rect 472636 4214 472664 69838
rect 474752 16574 474780 69906
rect 492680 68876 492732 68882
rect 492680 68818 492732 68824
rect 481640 68672 481692 68678
rect 481640 68614 481692 68620
rect 474752 16546 475792 16574
rect 473452 9036 473504 9042
rect 473452 8978 473504 8984
rect 472624 4208 472676 4214
rect 472624 4150 472676 4156
rect 472256 4072 472308 4078
rect 472256 4014 472308 4020
rect 472268 480 472296 4014
rect 473464 480 473492 8978
rect 474556 4208 474608 4214
rect 474556 4150 474608 4156
rect 474568 480 474596 4150
rect 475764 480 475792 16546
rect 478144 14544 478196 14550
rect 478144 14486 478196 14492
rect 476948 8968 477000 8974
rect 476948 8910 477000 8916
rect 476960 480 476988 8910
rect 478156 480 478184 14486
rect 480536 7880 480588 7886
rect 480536 7822 480588 7828
rect 479340 4004 479392 4010
rect 479340 3946 479392 3952
rect 479352 480 479380 3946
rect 480548 480 480576 7822
rect 481652 6914 481680 68614
rect 488540 68604 488592 68610
rect 488540 68546 488592 68552
rect 483020 68468 483072 68474
rect 483020 68410 483072 68416
rect 481732 17264 481784 17270
rect 481732 17206 481784 17212
rect 481744 16574 481772 17206
rect 483032 16574 483060 68410
rect 484400 67176 484452 67182
rect 484400 67118 484452 67124
rect 484412 16574 484440 67118
rect 485780 64388 485832 64394
rect 485780 64330 485832 64336
rect 485792 16574 485820 64330
rect 488552 16574 488580 68546
rect 489920 66972 489972 66978
rect 489920 66914 489972 66920
rect 481744 16546 482876 16574
rect 483032 16546 484072 16574
rect 484412 16546 485268 16574
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 482848 480 482876 16546
rect 484044 480 484072 16546
rect 485240 480 485268 16546
rect 486436 480 486464 16546
rect 487620 7336 487672 7342
rect 487620 7278 487672 7284
rect 487632 480 487660 7278
rect 488828 480 488856 16546
rect 489932 3398 489960 66914
rect 492692 16574 492720 68818
rect 503720 68808 503772 68814
rect 503720 68750 503772 68756
rect 500960 68400 501012 68406
rect 500960 68342 501012 68348
rect 496820 67312 496872 67318
rect 496820 67254 496872 67260
rect 496832 16574 496860 67254
rect 499580 18624 499632 18630
rect 499580 18566 499632 18572
rect 499592 16574 499620 18566
rect 500972 16574 501000 68342
rect 503732 16574 503760 68750
rect 528560 68740 528612 68746
rect 528560 68682 528612 68688
rect 506480 67244 506532 67250
rect 506480 67186 506532 67192
rect 492692 16546 493548 16574
rect 496832 16546 497136 16574
rect 499592 16546 500632 16574
rect 500972 16546 501828 16574
rect 503732 16546 504220 16574
rect 490012 10872 490064 10878
rect 490012 10814 490064 10820
rect 489920 3392 489972 3398
rect 489920 3334 489972 3340
rect 490024 1578 490052 10814
rect 492312 7676 492364 7682
rect 492312 7618 492364 7624
rect 491116 3392 491168 3398
rect 491116 3334 491168 3340
rect 489932 1550 490052 1578
rect 489932 480 489960 1550
rect 491128 480 491156 3334
rect 492324 480 492352 7618
rect 493520 480 493548 16546
rect 494704 13116 494756 13122
rect 494704 13058 494756 13064
rect 494716 480 494744 13058
rect 495900 7812 495952 7818
rect 495900 7754 495952 7760
rect 495912 480 495940 7754
rect 497108 480 497136 16546
rect 499396 11892 499448 11898
rect 499396 11834 499448 11840
rect 498200 11756 498252 11762
rect 498200 11698 498252 11704
rect 498212 480 498240 11698
rect 499408 480 499436 11834
rect 500604 480 500632 16546
rect 501800 480 501828 16546
rect 502984 5704 503036 5710
rect 502984 5646 503036 5652
rect 502996 480 503024 5646
rect 504192 480 504220 16546
rect 505376 7744 505428 7750
rect 505376 7686 505428 7692
rect 505388 480 505416 7686
rect 506492 3398 506520 67186
rect 507860 66904 507912 66910
rect 507860 66846 507912 66852
rect 507872 16574 507900 66846
rect 510620 65884 510672 65890
rect 510620 65826 510672 65832
rect 510632 16574 510660 65826
rect 524420 65816 524472 65822
rect 524420 65758 524472 65764
rect 517520 64320 517572 64326
rect 517520 64262 517572 64268
rect 514760 58676 514812 58682
rect 514760 58618 514812 58624
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 506572 5772 506624 5778
rect 506572 5714 506624 5720
rect 506480 3392 506532 3398
rect 506480 3334 506532 3340
rect 506584 2938 506612 5714
rect 507676 3392 507728 3398
rect 507676 3334 507728 3340
rect 506492 2910 506612 2938
rect 506492 480 506520 2910
rect 507688 480 507716 3334
rect 508884 480 508912 16546
rect 510068 5840 510120 5846
rect 510068 5782 510120 5788
rect 510080 480 510108 5782
rect 511276 480 511304 16546
rect 513564 5908 513616 5914
rect 513564 5850 513616 5856
rect 512460 4344 512512 4350
rect 512460 4286 512512 4292
rect 512472 480 512500 4286
rect 513576 480 513604 5850
rect 514772 480 514800 58618
rect 517532 16574 517560 64262
rect 521660 21412 521712 21418
rect 521660 21354 521712 21360
rect 521672 16574 521700 21354
rect 524432 16574 524460 65758
rect 528572 16574 528600 68682
rect 579620 68332 579672 68338
rect 579620 68274 579672 68280
rect 575480 65544 575532 65550
rect 575480 65486 575532 65492
rect 539600 64252 539652 64258
rect 539600 64194 539652 64200
rect 530584 62892 530636 62898
rect 530584 62834 530636 62840
rect 517532 16546 518388 16574
rect 521672 16546 521884 16574
rect 524432 16546 525472 16574
rect 528572 16546 529060 16574
rect 517152 5976 517204 5982
rect 517152 5918 517204 5924
rect 515956 4412 516008 4418
rect 515956 4354 516008 4360
rect 515968 480 515996 4354
rect 517164 480 517192 5918
rect 518360 480 518388 16546
rect 520740 6044 520792 6050
rect 520740 5986 520792 5992
rect 519544 4480 519596 4486
rect 519544 4422 519596 4428
rect 519556 480 519584 4422
rect 520752 480 520780 5986
rect 521856 480 521884 16546
rect 524236 6112 524288 6118
rect 524236 6054 524288 6060
rect 523040 4548 523092 4554
rect 523040 4490 523092 4496
rect 523052 480 523080 4490
rect 524248 480 524276 6054
rect 525444 480 525472 16546
rect 527824 6860 527876 6866
rect 527824 6802 527876 6808
rect 526628 4616 526680 4622
rect 526628 4558 526680 4564
rect 526640 480 526668 4558
rect 527836 480 527864 6802
rect 529032 480 529060 16546
rect 530124 4684 530176 4690
rect 530124 4626 530176 4632
rect 530136 480 530164 4626
rect 530596 3398 530624 62834
rect 535460 22772 535512 22778
rect 535460 22714 535512 22720
rect 535472 16574 535500 22714
rect 535472 16546 536144 16574
rect 531320 6792 531372 6798
rect 531320 6734 531372 6740
rect 530584 3392 530636 3398
rect 530584 3334 530636 3340
rect 531332 480 531360 6734
rect 534908 6724 534960 6730
rect 534908 6666 534960 6672
rect 533712 4752 533764 4758
rect 533712 4694 533764 4700
rect 532516 3392 532568 3398
rect 532516 3334 532568 3340
rect 532528 480 532556 3334
rect 533724 480 533752 4694
rect 534920 480 534948 6666
rect 536116 480 536144 16546
rect 538404 6656 538456 6662
rect 538404 6598 538456 6604
rect 537208 5500 537260 5506
rect 537208 5442 537260 5448
rect 537220 480 537248 5442
rect 538416 480 538444 6598
rect 539612 480 539640 64194
rect 546500 62824 546552 62830
rect 546500 62766 546552 62772
rect 542360 50380 542412 50386
rect 542360 50322 542412 50328
rect 542372 16574 542400 50322
rect 546512 16574 546540 62766
rect 575492 16574 575520 65486
rect 579632 16574 579660 68274
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 579894 33144 579950 33153
rect 579894 33079 579896 33088
rect 579948 33079 579950 33088
rect 579896 33050 579948 33056
rect 579896 20664 579948 20670
rect 579896 20606 579948 20612
rect 579908 19825 579936 20606
rect 579894 19816 579950 19825
rect 579894 19751 579950 19760
rect 542372 16546 543228 16574
rect 546512 16546 546724 16574
rect 575492 16546 576348 16574
rect 579632 16546 579844 16574
rect 541992 6588 542044 6594
rect 541992 6530 542044 6536
rect 540796 5432 540848 5438
rect 540796 5374 540848 5380
rect 540808 480 540836 5374
rect 542004 480 542032 6530
rect 543200 480 543228 16546
rect 545488 6520 545540 6526
rect 545488 6462 545540 6468
rect 544384 5364 544436 5370
rect 544384 5306 544436 5312
rect 544396 480 544424 5306
rect 545500 480 545528 6462
rect 546696 480 546724 16546
rect 563244 9648 563296 9654
rect 563244 9590 563296 9596
rect 549076 6452 549128 6458
rect 549076 6394 549128 6400
rect 547880 5296 547932 5302
rect 547880 5238 547932 5244
rect 547892 480 547920 5238
rect 549088 480 549116 6394
rect 552664 6384 552716 6390
rect 552664 6326 552716 6332
rect 551468 5228 551520 5234
rect 551468 5170 551520 5176
rect 550272 3936 550324 3942
rect 550272 3878 550324 3884
rect 550284 480 550312 3878
rect 551480 480 551508 5170
rect 552676 480 552704 6326
rect 556160 6316 556212 6322
rect 556160 6258 556212 6264
rect 554964 5160 555016 5166
rect 554964 5102 555016 5108
rect 553768 3868 553820 3874
rect 553768 3810 553820 3816
rect 553780 480 553808 3810
rect 554976 480 555004 5102
rect 556172 480 556200 6258
rect 559748 6248 559800 6254
rect 559748 6190 559800 6196
rect 558552 5092 558604 5098
rect 558552 5034 558604 5040
rect 557356 3800 557408 3806
rect 557356 3742 557408 3748
rect 557368 480 557396 3742
rect 558564 480 558592 5034
rect 559760 480 559788 6190
rect 562048 5024 562100 5030
rect 562048 4966 562100 4972
rect 560852 3732 560904 3738
rect 560852 3674 560904 3680
rect 560864 480 560892 3674
rect 562060 480 562088 4966
rect 563256 480 563284 9590
rect 570328 9512 570380 9518
rect 570328 9454 570380 9460
rect 566832 6180 566884 6186
rect 566832 6122 566884 6128
rect 565636 4956 565688 4962
rect 565636 4898 565688 4904
rect 564440 3664 564492 3670
rect 564440 3606 564492 3612
rect 564452 480 564480 3606
rect 565648 480 565676 4898
rect 566844 480 566872 6122
rect 569132 4888 569184 4894
rect 569132 4830 569184 4836
rect 568028 3596 568080 3602
rect 568028 3538 568080 3544
rect 568040 480 568068 3538
rect 569144 480 569172 4830
rect 570340 480 570368 9454
rect 573916 9308 573968 9314
rect 573916 9250 573968 9256
rect 572720 4820 572772 4826
rect 572720 4762 572772 4768
rect 571524 3528 571576 3534
rect 571524 3470 571576 3476
rect 571536 480 571564 3470
rect 572732 480 572760 4762
rect 573928 480 573956 9250
rect 575112 3460 575164 3466
rect 575112 3402 575164 3408
rect 575124 480 575152 3402
rect 576320 480 576348 16546
rect 577412 9240 577464 9246
rect 577412 9182 577464 9188
rect 577424 480 577452 9182
rect 578606 3632 578662 3641
rect 578606 3567 578662 3576
rect 578620 480 578648 3567
rect 579816 480 579844 16546
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 580184 5642 580212 6559
rect 580172 5636 580224 5642
rect 580172 5578 580224 5584
rect 582194 3768 582250 3777
rect 582194 3703 582250 3712
rect 580998 3496 581054 3505
rect 580998 3431 581054 3440
rect 581012 480 581040 3431
rect 582208 480 582236 3703
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
=======
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 100036 462 100340 490
rect 101048 480 101076 5170
rect 102244 480 102272 16546
rect 103440 6914 103468 70042
rect 103992 69086 104020 71726
rect 104164 69896 104216 69902
rect 104164 69838 104216 69844
rect 103980 69080 104032 69086
rect 103980 69022 104032 69028
rect 104176 14142 104204 69838
rect 104164 14136 104216 14142
rect 104164 14078 104216 14084
rect 104532 8968 104584 8974
rect 104532 8910 104584 8916
rect 103348 6886 103468 6914
rect 103348 480 103376 6886
rect 104544 480 104572 8910
rect 104728 5574 104756 71726
rect 105372 69086 105400 71726
rect 104808 69080 104860 69086
rect 104808 69022 104860 69028
rect 105360 69080 105412 69086
rect 105360 69022 105412 69028
rect 106096 69080 106148 69086
rect 106096 69022 106148 69028
rect 104716 5568 104768 5574
rect 104716 5510 104768 5516
rect 104820 4214 104848 69022
rect 105728 14136 105780 14142
rect 105728 14078 105780 14084
rect 104808 4208 104860 4214
rect 104808 4150 104860 4156
rect 105740 480 105768 14078
rect 106108 7614 106136 69022
rect 106096 7608 106148 7614
rect 106096 7550 106148 7556
rect 106200 4962 106228 71726
rect 106752 70174 106780 71726
rect 107396 71726 107464 71754
rect 107672 71862 108162 71890
rect 106740 70168 106792 70174
rect 106740 70110 106792 70116
rect 107396 66910 107424 71726
rect 107476 70100 107528 70106
rect 107476 70042 107528 70048
rect 107384 66904 107436 66910
rect 107384 66846 107436 66852
rect 107488 64874 107516 70042
rect 107568 69964 107620 69970
rect 107568 69906 107620 69912
rect 107580 69714 107608 69906
rect 107672 69834 107700 71862
rect 108832 71754 108860 72012
rect 107764 71726 108860 71754
rect 109132 71800 109184 71806
rect 109530 71754 109558 72012
rect 110228 71806 110256 72012
rect 109132 71742 109184 71748
rect 107660 69828 107712 69834
rect 107660 69770 107712 69776
rect 107580 69686 107700 69714
rect 107488 64846 107608 64874
rect 106188 4956 106240 4962
rect 106188 4898 106240 4904
rect 107580 3534 107608 64846
rect 107672 6914 107700 69686
rect 107764 16574 107792 71726
rect 107764 16546 107884 16574
rect 107672 6886 107792 6914
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 106936 480 106964 3470
rect 107764 3346 107792 6886
rect 107856 3466 107884 16546
rect 109144 3602 109172 71742
rect 109236 71726 109558 71754
rect 110216 71800 110268 71806
rect 110925 71754 110953 72012
rect 111623 71754 111651 72012
rect 112321 71754 112349 72012
rect 113019 71754 113047 72012
rect 113717 71754 113745 72012
rect 114414 71754 114442 72012
rect 110216 71742 110268 71748
rect 110524 71726 110953 71754
rect 110984 71726 111651 71754
rect 111904 71726 112349 71754
rect 112456 71726 113047 71754
rect 113284 71726 113745 71754
rect 114388 71726 114442 71754
rect 114560 71800 114612 71806
rect 114560 71742 114612 71748
rect 115112 71754 115140 72012
rect 115810 71806 115838 72012
rect 115798 71800 115850 71806
rect 109132 3596 109184 3602
rect 109132 3538 109184 3544
rect 109236 3534 109264 71726
rect 109316 4208 109368 4214
rect 109316 4150 109368 4156
rect 109224 3528 109276 3534
rect 109224 3470 109276 3476
rect 107844 3460 107896 3466
rect 107844 3402 107896 3408
rect 107764 3318 108160 3346
rect 108132 480 108160 3318
rect 109328 480 109356 4150
rect 110524 3670 110552 71726
rect 110984 64874 111012 71726
rect 111708 69828 111760 69834
rect 111708 69770 111760 69776
rect 110616 64846 111012 64874
rect 110616 3738 110644 64846
rect 111616 5092 111668 5098
rect 111616 5034 111668 5040
rect 110604 3732 110656 3738
rect 110604 3674 110656 3680
rect 110512 3664 110564 3670
rect 110512 3606 110564 3612
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 110524 480 110552 3470
rect 111628 480 111656 5034
rect 111720 3534 111748 69770
rect 111800 69284 111852 69290
rect 111800 69226 111852 69232
rect 111812 68338 111840 69226
rect 111800 68332 111852 68338
rect 111800 68274 111852 68280
rect 111904 3806 111932 71726
rect 112456 64874 112484 71726
rect 111996 64846 112484 64874
rect 111996 3874 112024 64846
rect 112812 5568 112864 5574
rect 112812 5510 112864 5516
rect 111984 3868 112036 3874
rect 111984 3810 112036 3816
rect 111892 3800 111944 3806
rect 111892 3742 111944 3748
rect 111708 3528 111760 3534
rect 111708 3470 111760 3476
rect 112824 480 112852 5510
rect 113284 3534 113312 71726
rect 114388 69290 114416 71726
rect 114468 69964 114520 69970
rect 114468 69906 114520 69912
rect 114376 69284 114428 69290
rect 114376 69226 114428 69232
rect 114480 3534 114508 69906
rect 113272 3528 113324 3534
rect 113272 3470 113324 3476
rect 114008 3528 114060 3534
rect 114008 3470 114060 3476
rect 114468 3528 114520 3534
rect 114468 3470 114520 3476
rect 114020 480 114048 3470
rect 114572 3466 114600 71742
rect 115112 71726 115152 71754
rect 115798 71742 115850 71748
rect 116032 71800 116084 71806
rect 116508 71754 116536 72012
rect 117206 71806 117234 72012
rect 116032 71742 116084 71748
rect 114652 65680 114704 65686
rect 114652 65622 114704 65628
rect 114664 16574 114692 65622
rect 115124 65550 115152 71726
rect 115112 65544 115164 65550
rect 115112 65486 115164 65492
rect 114664 16546 114784 16574
rect 114560 3460 114612 3466
rect 114560 3402 114612 3408
rect 114756 490 114784 16546
rect 116044 4146 116072 71742
rect 116136 71726 116536 71754
rect 117194 71800 117246 71806
rect 117194 71742 117246 71748
rect 117320 71800 117372 71806
rect 117903 71754 117931 72012
rect 118601 71806 118629 72012
rect 117320 71742 117372 71748
rect 116032 4140 116084 4146
rect 116032 4082 116084 4088
rect 116136 4078 116164 71726
rect 116400 7608 116452 7614
rect 116400 7550 116452 7556
rect 116124 4072 116176 4078
rect 116124 4014 116176 4020
rect 115032 598 115244 626
rect 115032 490 115060 598
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 462 115060 490
rect 115216 480 115244 598
rect 116412 480 116440 7550
rect 116492 4956 116544 4962
rect 116492 4898 116544 4904
rect 116504 2922 116532 4898
rect 117332 3330 117360 71742
rect 117424 71726 117931 71754
rect 118589 71800 118641 71806
rect 118589 71742 118641 71748
rect 118792 71800 118844 71806
rect 119299 71754 119327 72012
rect 119997 71806 120025 72012
rect 118792 71742 118844 71748
rect 117424 3398 117452 71726
rect 118804 6914 118832 71742
rect 118712 6886 118832 6914
rect 118988 71726 119327 71754
rect 119985 71800 120037 71806
rect 119985 71742 120037 71748
rect 120172 71800 120224 71806
rect 120695 71754 120723 72012
rect 121392 71806 121420 72012
rect 120172 71742 120224 71748
rect 117412 3392 117464 3398
rect 117412 3334 117464 3340
rect 117320 3324 117372 3330
rect 117320 3266 117372 3272
rect 118712 3194 118740 6886
rect 118792 4888 118844 4894
rect 118792 4830 118844 4836
rect 118700 3188 118752 3194
rect 118700 3130 118752 3136
rect 117596 3052 117648 3058
rect 117596 2994 117648 3000
rect 116492 2916 116544 2922
rect 116492 2858 116544 2864
rect 117608 480 117636 2994
rect 118804 480 118832 4830
rect 118988 3262 119016 71726
rect 119344 70236 119396 70242
rect 119344 70178 119396 70184
rect 118976 3256 119028 3262
rect 118976 3198 119028 3204
rect 119356 3058 119384 70178
rect 119344 3052 119396 3058
rect 119344 2994 119396 3000
rect 120184 2990 120212 71742
rect 120276 71726 120723 71754
rect 121380 71800 121432 71806
rect 122090 71754 122118 72012
rect 122788 71754 122816 72012
rect 123486 71754 123514 72012
rect 124184 71754 124212 72012
rect 124881 71754 124909 72012
rect 121380 71742 121432 71748
rect 121564 71726 122118 71754
rect 122208 71726 122816 71754
rect 122944 71726 123514 71754
rect 124140 71726 124212 71754
rect 124876 71726 124909 71754
rect 125579 71754 125607 72012
rect 126277 71754 126305 72012
rect 125579 71726 125640 71754
rect 120276 3126 120304 71726
rect 121368 70304 121420 70310
rect 121368 70246 121420 70252
rect 121380 6914 121408 70246
rect 121104 6886 121408 6914
rect 120264 3120 120316 3126
rect 120264 3062 120316 3068
rect 120172 2984 120224 2990
rect 120172 2926 120224 2932
rect 119896 2916 119948 2922
rect 119896 2858 119948 2864
rect 119908 480 119936 2858
rect 121104 480 121132 6886
rect 121564 3466 121592 71726
rect 122208 64874 122236 71726
rect 122840 70168 122892 70174
rect 122840 70110 122892 70116
rect 121656 64846 122236 64874
rect 121656 3534 121684 64846
rect 122288 4820 122340 4826
rect 122288 4762 122340 4768
rect 121644 3528 121696 3534
rect 121644 3470 121696 3476
rect 121552 3460 121604 3466
rect 121552 3402 121604 3408
rect 122300 480 122328 4762
rect 122852 626 122880 70110
rect 122944 2854 122972 71726
rect 124140 69902 124168 71726
rect 124876 70038 124904 71726
rect 125612 70106 125640 71726
rect 126256 71726 126305 71754
rect 126975 71754 127003 72012
rect 127673 71754 127701 72012
rect 126975 71726 127020 71754
rect 125600 70100 125652 70106
rect 125600 70042 125652 70048
rect 124864 70032 124916 70038
rect 124864 69974 124916 69980
rect 124128 69896 124180 69902
rect 124128 69838 124180 69844
rect 126256 69834 126284 71726
rect 126992 69970 127020 71726
rect 127636 71726 127701 71754
rect 128370 71754 128398 72012
rect 129068 71754 129096 72012
rect 128370 71726 128400 71754
rect 127636 70242 127664 71726
rect 128372 70310 128400 71726
rect 129016 71726 129096 71754
rect 129766 71754 129794 72012
rect 130464 71754 130492 72012
rect 131162 71754 131190 72012
rect 131859 71754 131887 72012
rect 129766 71726 129872 71754
rect 130464 71726 130516 71754
rect 128360 70304 128412 70310
rect 128360 70246 128412 70252
rect 127624 70236 127676 70242
rect 127624 70178 127676 70184
rect 126980 69964 127032 69970
rect 126980 69906 127032 69912
rect 126244 69828 126296 69834
rect 126244 69770 126296 69776
rect 126888 69420 126940 69426
rect 126888 69362 126940 69368
rect 125508 69080 125560 69086
rect 125508 69022 125560 69028
rect 125520 3534 125548 69022
rect 126900 3534 126928 69362
rect 129016 69086 129044 71726
rect 129648 69896 129700 69902
rect 129648 69838 129700 69844
rect 129004 69080 129056 69086
rect 129004 69022 129056 69028
rect 129556 9240 129608 9246
rect 129556 9182 129608 9188
rect 129568 3534 129596 9182
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 129556 3528 129608 3534
rect 129556 3470 129608 3476
rect 122932 2848 122984 2854
rect 122932 2790 122984 2796
rect 122852 598 123064 626
rect 123036 490 123064 598
rect 123312 598 123524 626
rect 123312 490 123340 598
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
<<<<<<< HEAD
=======
rect 123036 462 123340 490
rect 123496 480 123524 598
rect 124692 480 124720 3470
rect 125888 480 125916 3470
rect 126992 480 127020 3470
rect 128176 3460 128228 3466
rect 128176 3402 128228 3408
rect 128188 480 128216 3402
rect 129660 3346 129688 69838
rect 129844 3505 129872 71726
rect 130488 69766 130516 71726
rect 131132 71726 131190 71754
rect 131224 71726 131887 71754
rect 132557 71754 132585 72012
rect 133255 71754 133283 72012
rect 133953 71754 133981 72012
rect 134651 71754 134679 72012
rect 132557 71726 132632 71754
rect 131028 69828 131080 69834
rect 131028 69770 131080 69776
rect 130476 69760 130528 69766
rect 130476 69702 130528 69708
rect 131040 3534 131068 69770
rect 131132 3641 131160 71726
rect 131224 3777 131252 71726
rect 131764 3868 131816 3874
rect 131764 3810 131816 3816
rect 131210 3768 131266 3777
rect 131210 3703 131266 3712
rect 131118 3632 131174 3641
rect 131118 3567 131174 3576
rect 130568 3528 130620 3534
rect 129830 3496 129886 3505
rect 130568 3470 130620 3476
rect 131028 3528 131080 3534
rect 131028 3470 131080 3476
rect 129830 3431 129886 3440
rect 129384 3318 129688 3346
rect 129384 480 129412 3318
rect 130580 480 130608 3470
rect 131776 480 131804 3810
rect 132604 3369 132632 71726
rect 133248 71726 133283 71754
rect 133892 71726 133981 71754
rect 134628 71726 134679 71754
rect 135348 71754 135376 72012
rect 136046 71754 136074 72012
rect 135348 71726 135392 71754
rect 133248 69698 133276 71726
rect 133236 69692 133288 69698
rect 133236 69634 133288 69640
rect 133892 69426 133920 71726
rect 134628 69902 134656 71726
rect 135168 70032 135220 70038
rect 135168 69974 135220 69980
rect 134616 69896 134668 69902
rect 134616 69838 134668 69844
rect 133880 69420 133932 69426
rect 133880 69362 133932 69368
rect 133788 69080 133840 69086
rect 133788 69022 133840 69028
rect 133800 3534 133828 69022
rect 134524 68604 134576 68610
rect 134524 68546 134576 68552
rect 132960 3528 133012 3534
rect 132960 3470 133012 3476
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 132590 3360 132646 3369
rect 132590 3295 132646 3304
rect 132972 480 133000 3470
rect 134536 3466 134564 68546
rect 134524 3460 134576 3466
rect 134524 3402 134576 3408
rect 135180 3194 135208 69974
rect 135364 69086 135392 71726
rect 135456 71726 136074 71754
rect 135352 69080 135404 69086
rect 135352 69022 135404 69028
rect 135260 3800 135312 3806
rect 135260 3742 135312 3748
rect 134156 3188 134208 3194
rect 134156 3130 134208 3136
rect 135168 3188 135220 3194
rect 135168 3130 135220 3136
rect 134168 480 134196 3130
rect 135272 480 135300 3742
rect 135456 2922 135484 71726
rect 136744 69086 136772 72012
rect 137442 71754 137470 72012
rect 138140 71754 138168 72012
rect 137442 71726 137784 71754
rect 136732 69080 136784 69086
rect 136732 69022 136784 69028
rect 137756 3058 137784 71726
rect 138124 71726 138168 71754
rect 138837 71754 138865 72012
rect 139535 71754 139563 72012
rect 140233 71754 140261 72012
rect 140931 71754 140959 72012
rect 141629 71754 141657 72012
rect 142326 71754 142354 72012
rect 143024 71754 143052 72012
rect 143722 71754 143750 72012
rect 144420 71754 144448 72012
rect 145118 71754 145146 72012
rect 138837 71726 139256 71754
rect 139535 71726 139624 71754
rect 140233 71726 140636 71754
rect 140931 71726 141004 71754
rect 141629 71726 141924 71754
rect 142326 71726 142384 71754
rect 143024 71726 143396 71754
rect 143722 71726 143764 71754
rect 144420 71726 144776 71754
rect 137928 70168 137980 70174
rect 137928 70110 137980 70116
rect 137836 69080 137888 69086
rect 137836 69022 137888 69028
rect 137848 3398 137876 69022
rect 137836 3392 137888 3398
rect 137836 3334 137888 3340
rect 137744 3052 137796 3058
rect 137744 2994 137796 3000
rect 137940 2938 137968 70110
rect 138124 69086 138152 71726
rect 138112 69080 138164 69086
rect 138112 69022 138164 69028
rect 139228 3602 139256 71726
rect 139596 69086 139624 71726
rect 139308 69080 139360 69086
rect 139308 69022 139360 69028
rect 139584 69080 139636 69086
rect 139584 69022 139636 69028
rect 139216 3596 139268 3602
rect 139216 3538 139268 3544
rect 139320 3466 139348 69022
rect 140608 3942 140636 71726
rect 140976 69086 141004 71726
rect 140688 69080 140740 69086
rect 140688 69022 140740 69028
rect 140964 69080 141016 69086
rect 140964 69022 141016 69028
rect 140596 3936 140648 3942
rect 140596 3878 140648 3884
rect 140700 3670 140728 69022
rect 141896 6186 141924 71726
rect 141976 70304 142028 70310
rect 141976 70246 142028 70252
rect 141884 6180 141936 6186
rect 141884 6122 141936 6128
rect 140688 3664 140740 3670
rect 140688 3606 140740 3612
rect 141988 3534 142016 70246
rect 142356 69086 142384 71726
rect 142068 69080 142120 69086
rect 142068 69022 142120 69028
rect 142344 69080 142396 69086
rect 142344 69022 142396 69028
rect 142080 3738 142108 69022
rect 143368 4554 143396 71726
rect 143736 69086 143764 71726
rect 143448 69080 143500 69086
rect 143448 69022 143500 69028
rect 143724 69080 143776 69086
rect 143724 69022 143776 69028
rect 144644 69080 144696 69086
rect 144644 69022 144696 69028
rect 143356 4548 143408 4554
rect 143356 4490 143408 4496
rect 143460 4486 143488 69022
rect 144656 16574 144684 69022
rect 144564 16546 144684 16574
rect 144564 4622 144592 16546
rect 144748 11778 144776 71726
rect 145116 71726 145146 71754
rect 145815 71754 145843 72012
rect 146513 71754 146541 72012
rect 145815 71726 146248 71754
rect 144828 70236 144880 70242
rect 144828 70178 144880 70184
rect 144656 11750 144776 11778
rect 144656 4690 144684 11750
rect 144840 6914 144868 70178
rect 145116 69086 145144 71726
rect 145104 69080 145156 69086
rect 145104 69022 145156 69028
rect 146116 69080 146168 69086
rect 146116 69022 146168 69028
rect 144748 6886 144868 6914
rect 144644 4684 144696 4690
rect 144644 4626 144696 4632
rect 144552 4616 144604 4622
rect 144552 4558 144604 4564
rect 143448 4480 143500 4486
rect 143448 4422 143500 4428
rect 142068 3732 142120 3738
rect 142068 3674 142120 3680
rect 141240 3528 141292 3534
rect 141240 3470 141292 3476
rect 141976 3528 142028 3534
rect 141976 3470 142028 3476
rect 142434 3496 142490 3505
rect 139308 3460 139360 3466
rect 139308 3402 139360 3408
rect 140044 3392 140096 3398
rect 138846 3360 138902 3369
rect 140044 3334 140096 3340
rect 138846 3295 138902 3304
rect 135444 2916 135496 2922
rect 135444 2858 135496 2864
rect 136456 2916 136508 2922
rect 136456 2858 136508 2864
rect 137664 2910 137968 2938
rect 136468 480 136496 2858
rect 137664 480 137692 2910
rect 138860 480 138888 3295
rect 140056 480 140084 3334
rect 141252 480 141280 3470
rect 142434 3431 142490 3440
rect 142448 480 142476 3431
rect 143540 3052 143592 3058
rect 143540 2994 143592 3000
rect 143552 480 143580 2994
rect 144748 480 144776 6886
rect 146128 4758 146156 69022
rect 146220 5506 146248 71726
rect 146496 71726 146541 71754
rect 147211 71754 147239 72012
rect 147909 71754 147937 72012
rect 148607 71754 148635 72012
rect 149304 71754 149332 72012
rect 150002 71754 150030 72012
rect 150700 71754 150728 72012
rect 151398 71754 151426 72012
rect 152096 71754 152124 72012
rect 152793 71754 152821 72012
rect 153491 71754 153519 72012
rect 147211 71726 147536 71754
rect 147909 71726 147996 71754
rect 148607 71726 148824 71754
rect 149304 71726 149376 71754
rect 150002 71726 150388 71754
rect 150700 71726 150756 71754
rect 151398 71726 151676 71754
rect 152096 71726 152136 71754
rect 152793 71726 153148 71754
rect 146496 69086 146524 71726
rect 146484 69080 146536 69086
rect 146484 69022 146536 69028
rect 146208 5500 146260 5506
rect 146208 5442 146260 5448
rect 147508 5370 147536 71726
rect 147968 69086 147996 71726
rect 147588 69080 147640 69086
rect 147588 69022 147640 69028
rect 147956 69080 148008 69086
rect 147956 69022 148008 69028
rect 147600 5438 147628 69022
rect 147588 5432 147640 5438
rect 147588 5374 147640 5380
rect 147496 5364 147548 5370
rect 147496 5306 147548 5312
rect 148796 5234 148824 71726
rect 148968 70372 149020 70378
rect 148968 70314 149020 70320
rect 148876 69080 148928 69086
rect 148876 69022 148928 69028
rect 148888 5302 148916 69022
rect 148876 5296 148928 5302
rect 148876 5238 148928 5244
rect 148784 5228 148836 5234
rect 148784 5170 148836 5176
rect 146116 4752 146168 4758
rect 146116 4694 146168 4700
rect 148980 3534 149008 70314
rect 149348 69086 149376 71726
rect 149336 69080 149388 69086
rect 149336 69022 149388 69028
rect 150256 69080 150308 69086
rect 150256 69022 150308 69028
rect 150268 5166 150296 69022
rect 150256 5160 150308 5166
rect 150256 5102 150308 5108
rect 150360 5098 150388 71726
rect 150728 69086 150756 71726
rect 150716 69080 150768 69086
rect 150716 69022 150768 69028
rect 150348 5092 150400 5098
rect 150348 5034 150400 5040
rect 151648 4962 151676 71726
rect 152108 69086 152136 71726
rect 151728 69080 151780 69086
rect 151728 69022 151780 69028
rect 152096 69080 152148 69086
rect 152096 69022 152148 69028
rect 153016 69080 153068 69086
rect 153016 69022 153068 69028
rect 151740 5030 151768 69022
rect 151728 5024 151780 5030
rect 151728 4966 151780 4972
rect 151636 4956 151688 4962
rect 151636 4898 151688 4904
rect 153028 4894 153056 69022
rect 153016 4888 153068 4894
rect 153016 4830 153068 4836
rect 153120 4826 153148 71726
rect 153488 71726 153519 71754
rect 154189 71754 154217 72012
rect 154887 71754 154915 72012
rect 154189 71726 154252 71754
rect 153488 69086 153516 71726
rect 154224 69766 154252 71726
rect 154868 71726 154915 71754
rect 155585 71754 155613 72012
rect 156282 71754 156310 72012
rect 156980 71754 157008 72012
rect 157678 71754 157706 72012
rect 158376 71754 158404 72012
rect 159074 71754 159102 72012
rect 159771 71754 159799 72012
rect 160469 71754 160497 72012
rect 161167 71754 161195 72012
rect 161865 71754 161893 72012
rect 155585 71726 155816 71754
rect 156282 71726 156368 71754
rect 156980 71726 157288 71754
rect 157678 71726 157748 71754
rect 158376 71726 158668 71754
rect 159074 71726 159128 71754
rect 159771 71726 160048 71754
rect 160469 71726 160508 71754
rect 161167 71726 161336 71754
rect 154212 69760 154264 69766
rect 154212 69702 154264 69708
rect 154868 69426 154896 71726
rect 154856 69420 154908 69426
rect 154856 69362 154908 69368
rect 153476 69080 153528 69086
rect 153476 69022 153528 69028
rect 154488 69080 154540 69086
rect 154488 69022 154540 69028
rect 153108 4820 153160 4826
rect 153108 4762 153160 4768
rect 154500 4282 154528 69022
rect 155788 6662 155816 71726
rect 155868 69624 155920 69630
rect 155868 69566 155920 69572
rect 155776 6656 155828 6662
rect 155776 6598 155828 6604
rect 154488 4276 154540 4282
rect 154488 4218 154540 4224
rect 154212 3664 154264 3670
rect 154212 3606 154264 3612
rect 150624 3596 150676 3602
rect 150624 3538 150676 3544
rect 153016 3596 153068 3602
rect 153016 3538 153068 3544
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 145932 3460 145984 3466
rect 145932 3402 145984 3408
rect 145944 480 145972 3402
rect 147128 3392 147180 3398
rect 147128 3334 147180 3340
rect 147140 480 147168 3334
rect 148336 480 148364 3470
rect 149532 480 149560 3470
rect 150636 480 150664 3538
rect 151820 2984 151872 2990
rect 151820 2926 151872 2932
rect 151832 480 151860 2926
rect 153028 480 153056 3538
rect 154224 480 154252 3606
rect 155880 3398 155908 69566
rect 156340 69358 156368 71726
rect 156328 69352 156380 69358
rect 156328 69294 156380 69300
rect 157260 6594 157288 71726
rect 157720 69562 157748 71726
rect 157708 69556 157760 69562
rect 157708 69498 157760 69504
rect 158640 10606 158668 71726
rect 159100 69086 159128 71726
rect 159088 69080 159140 69086
rect 159088 69022 159140 69028
rect 159916 69080 159968 69086
rect 159916 69022 159968 69028
rect 158628 10600 158680 10606
rect 158628 10542 158680 10548
rect 159928 10538 159956 69022
rect 159916 10532 159968 10538
rect 159916 10474 159968 10480
rect 157248 6588 157300 6594
rect 157248 6530 157300 6536
rect 160020 6526 160048 71726
rect 160480 69086 160508 71726
rect 160468 69080 160520 69086
rect 160468 69022 160520 69028
rect 160744 12096 160796 12102
rect 160744 12038 160796 12044
rect 160008 6520 160060 6526
rect 160008 6462 160060 6468
rect 157800 3936 157852 3942
rect 157800 3878 157852 3884
rect 158904 3936 158956 3942
rect 158904 3878 158956 3884
rect 156604 3664 156656 3670
rect 156604 3606 156656 3612
rect 155408 3392 155460 3398
rect 155408 3334 155460 3340
rect 155868 3392 155920 3398
rect 155868 3334 155920 3340
rect 155420 480 155448 3334
rect 156616 480 156644 3606
rect 157812 480 157840 3878
rect 158916 480 158944 3878
rect 160100 3732 160152 3738
rect 160100 3674 160152 3680
rect 160112 480 160140 3674
rect 160756 2990 160784 12038
rect 161308 10402 161336 71726
rect 161860 71726 161893 71754
rect 162563 71754 162591 72012
rect 163260 71754 163288 72012
rect 162563 71726 162808 71754
rect 161860 69086 161888 71726
rect 161388 69080 161440 69086
rect 161388 69022 161440 69028
rect 161848 69080 161900 69086
rect 161848 69022 161900 69028
rect 162676 69080 162728 69086
rect 162676 69022 162728 69028
rect 161400 10470 161428 69022
rect 162124 18624 162176 18630
rect 162124 18566 162176 18572
rect 161388 10464 161440 10470
rect 161388 10406 161440 10412
rect 161296 10396 161348 10402
rect 161296 10338 161348 10344
rect 162136 3874 162164 18566
rect 162688 12034 162716 69022
rect 162676 12028 162728 12034
rect 162676 11970 162728 11976
rect 162492 10668 162544 10674
rect 162492 10610 162544 10616
rect 162124 3868 162176 3874
rect 162124 3810 162176 3816
rect 161296 3392 161348 3398
rect 161296 3334 161348 3340
rect 160744 2984 160796 2990
rect 160744 2926 160796 2932
rect 161308 480 161336 3334
rect 162504 480 162532 10610
rect 162780 10334 162808 71726
rect 163240 71726 163288 71754
rect 163958 71754 163986 72012
rect 164656 71754 164684 72012
rect 165354 71754 165382 72012
rect 166052 71754 166080 72012
rect 166749 71754 166777 72012
rect 167447 71754 167475 72012
rect 168145 71754 168173 72012
rect 168843 71754 168871 72012
rect 169541 71754 169569 72012
rect 170238 71754 170266 72012
rect 163958 71726 164004 71754
rect 164656 71726 164740 71754
rect 165354 71726 165568 71754
rect 166052 71726 166120 71754
rect 166749 71726 166948 71754
rect 167447 71726 167500 71754
rect 168145 71726 168236 71754
rect 168843 71726 168880 71754
rect 169541 71726 169616 71754
rect 163240 69290 163268 71726
rect 163976 70106 164004 71726
rect 163964 70100 164016 70106
rect 163964 70042 164016 70048
rect 164712 69494 164740 71726
rect 164700 69488 164752 69494
rect 164700 69430 164752 69436
rect 163228 69284 163280 69290
rect 163228 69226 163280 69232
rect 164148 15972 164200 15978
rect 164148 15914 164200 15920
rect 162768 10328 162820 10334
rect 162768 10270 162820 10276
rect 164160 3398 164188 15914
rect 165540 11898 165568 71726
rect 166092 69086 166120 71726
rect 166080 69080 166132 69086
rect 166080 69022 166132 69028
rect 166816 69080 166868 69086
rect 166816 69022 166868 69028
rect 165528 11892 165580 11898
rect 165528 11834 165580 11840
rect 166828 6390 166856 69022
rect 166816 6384 166868 6390
rect 166816 6326 166868 6332
rect 166920 6322 166948 71726
rect 167472 69086 167500 71726
rect 167460 69080 167512 69086
rect 167460 69022 167512 69028
rect 167184 6452 167236 6458
rect 167184 6394 167236 6400
rect 166908 6316 166960 6322
rect 166908 6258 166960 6264
rect 164884 6180 164936 6186
rect 164884 6122 164936 6128
rect 163688 3392 163740 3398
rect 163688 3334 163740 3340
rect 164148 3392 164200 3398
rect 164148 3334 164200 3340
rect 163700 480 163728 3334
rect 164896 480 164924 6122
rect 166080 3188 166132 3194
rect 166080 3130 166132 3136
rect 166092 480 166120 3130
rect 167196 480 167224 6394
rect 168208 6186 168236 71726
rect 168852 69086 168880 71726
rect 168288 69080 168340 69086
rect 168288 69022 168340 69028
rect 168840 69080 168892 69086
rect 168840 69022 168892 69028
rect 168300 6254 168328 69022
rect 169588 13530 169616 71726
rect 170232 71726 170266 71754
rect 170936 71754 170964 72012
rect 171634 71754 171662 72012
rect 170936 71726 171088 71754
rect 170232 69086 170260 71726
rect 169668 69080 169720 69086
rect 169668 69022 169720 69028
rect 170220 69080 170272 69086
rect 170220 69022 170272 69028
rect 170956 69080 171008 69086
rect 170956 69022 171008 69028
rect 169576 13524 169628 13530
rect 169576 13466 169628 13472
rect 169680 12306 169708 69022
rect 170968 14754 170996 69022
rect 170956 14748 171008 14754
rect 170956 14690 171008 14696
rect 170404 14544 170456 14550
rect 170404 14486 170456 14492
rect 169668 12300 169720 12306
rect 169668 12242 169720 12248
rect 169576 12164 169628 12170
rect 169576 12106 169628 12112
rect 168288 6248 168340 6254
rect 168288 6190 168340 6196
rect 168196 6180 168248 6186
rect 168196 6122 168248 6128
rect 168380 4480 168432 4486
rect 168380 4422 168432 4428
rect 168392 480 168420 4422
rect 169588 480 169616 12106
rect 170416 3194 170444 14486
rect 171060 12238 171088 71726
rect 171612 71726 171662 71754
rect 172332 71754 172360 72012
rect 173030 71754 173058 72012
rect 173727 71754 173755 72012
rect 174425 71754 174453 72012
rect 175123 71754 175151 72012
rect 175821 71754 175849 72012
rect 176519 71754 176547 72012
rect 177216 71754 177244 72012
rect 177914 71754 177942 72012
rect 178612 71754 178640 72012
rect 172332 71726 172376 71754
rect 173030 71726 173112 71754
rect 173727 71726 173756 71754
rect 174425 71726 174492 71754
rect 175123 71726 175228 71754
rect 175821 71726 175872 71754
rect 176519 71726 176608 71754
rect 177216 71726 177252 71754
rect 171612 69086 171640 71726
rect 171600 69080 171652 69086
rect 171600 69022 171652 69028
rect 172348 68814 172376 71726
rect 173084 69154 173112 71726
rect 173072 69148 173124 69154
rect 173072 69090 173124 69096
rect 173164 69080 173216 69086
rect 173164 69022 173216 69028
rect 172336 68808 172388 68814
rect 172336 68750 172388 68756
rect 173176 16046 173204 69022
rect 173256 16108 173308 16114
rect 173256 16050 173308 16056
rect 173164 16040 173216 16046
rect 173164 15982 173216 15988
rect 171048 12232 171100 12238
rect 171048 12174 171100 12180
rect 171968 4548 172020 4554
rect 171968 4490 172020 4496
rect 170772 3868 170824 3874
rect 170772 3810 170824 3816
rect 170404 3188 170456 3194
rect 170404 3130 170456 3136
rect 170784 480 170812 3810
rect 171980 480 172008 4490
rect 173268 3806 173296 16050
rect 173624 13728 173676 13734
rect 173624 13670 173676 13676
rect 173256 3800 173308 3806
rect 173256 3742 173308 3748
rect 173636 3398 173664 13670
rect 173728 13394 173756 71726
rect 173808 69148 173860 69154
rect 173808 69090 173860 69096
rect 173820 13462 173848 69090
rect 174464 69086 174492 71726
rect 174452 69080 174504 69086
rect 174452 69022 174504 69028
rect 175096 69080 175148 69086
rect 175096 69022 175148 69028
rect 175108 47598 175136 69022
rect 175096 47592 175148 47598
rect 175096 47534 175148 47540
rect 175096 17264 175148 17270
rect 175096 17206 175148 17212
rect 173808 13456 173860 13462
rect 173808 13398 173860 13404
rect 173716 13388 173768 13394
rect 173716 13330 173768 13336
rect 175108 3398 175136 17206
rect 175200 14686 175228 71726
rect 175844 69086 175872 71726
rect 175832 69080 175884 69086
rect 175832 69022 175884 69028
rect 176476 69080 176528 69086
rect 176476 69022 176528 69028
rect 176488 49026 176516 69022
rect 176476 49020 176528 49026
rect 176476 48962 176528 48968
rect 175188 14680 175240 14686
rect 175188 14622 175240 14628
rect 176580 11966 176608 71726
rect 177224 68746 177252 71726
rect 177776 71726 177942 71754
rect 178604 71726 178640 71754
rect 179310 71754 179338 72012
rect 180008 71754 180036 72012
rect 179310 71726 179368 71754
rect 177212 68740 177264 68746
rect 177212 68682 177264 68688
rect 177304 68536 177356 68542
rect 177304 68478 177356 68484
rect 176568 11960 176620 11966
rect 176568 11902 176620 11908
rect 175464 4616 175516 4622
rect 175464 4558 175516 4564
rect 173164 3392 173216 3398
rect 173164 3334 173216 3340
rect 173624 3392 173676 3398
rect 173624 3334 173676 3340
rect 174268 3392 174320 3398
rect 174268 3334 174320 3340
rect 175096 3392 175148 3398
rect 175096 3334 175148 3340
rect 173176 480 173204 3334
rect 174280 480 174308 3334
rect 175476 480 175504 4558
rect 177316 3942 177344 68478
rect 177776 13326 177804 71726
rect 178604 69086 178632 71726
rect 178592 69080 178644 69086
rect 178592 69022 178644 69028
rect 179236 69080 179288 69086
rect 179236 69022 179288 69028
rect 177856 17468 177908 17474
rect 177856 17410 177908 17416
rect 177764 13320 177816 13326
rect 177764 13262 177816 13268
rect 177304 3936 177356 3942
rect 177304 3878 177356 3884
rect 177868 3398 177896 17410
rect 178684 17332 178736 17338
rect 178684 17274 178736 17280
rect 178696 3874 178724 17274
rect 179248 14618 179276 69022
rect 179236 14612 179288 14618
rect 179236 14554 179288 14560
rect 179340 7070 179368 71726
rect 179984 71726 180036 71754
rect 180705 71754 180733 72012
rect 181403 71754 181431 72012
rect 182101 71754 182129 72012
rect 180705 71726 180748 71754
rect 181403 71726 181484 71754
rect 179984 69086 180012 71726
rect 179972 69080 180024 69086
rect 179972 69022 180024 69028
rect 180616 69080 180668 69086
rect 180616 69022 180668 69028
rect 180248 9512 180300 9518
rect 180248 9454 180300 9460
rect 179328 7064 179380 7070
rect 179328 7006 179380 7012
rect 179052 4684 179104 4690
rect 179052 4626 179104 4632
rect 178684 3868 178736 3874
rect 178684 3810 178736 3816
rect 177948 3800 178000 3806
rect 177948 3742 178000 3748
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 177856 3392 177908 3398
rect 177856 3334 177908 3340
rect 176672 480 176700 3334
rect 177960 1986 177988 3742
rect 177868 1958 177988 1986
rect 177868 480 177896 1958
rect 179064 480 179092 4626
rect 180260 480 180288 9454
rect 180628 7138 180656 69022
rect 180720 7206 180748 71726
rect 181456 69086 181484 71726
rect 182008 71726 182129 71754
rect 182799 71754 182827 72012
rect 183497 71754 183525 72012
rect 182799 71726 182864 71754
rect 181444 69080 181496 69086
rect 181444 69022 181496 69028
rect 181904 12368 181956 12374
rect 181904 12310 181956 12316
rect 180708 7200 180760 7206
rect 180708 7142 180760 7148
rect 180616 7132 180668 7138
rect 180616 7074 180668 7080
rect 181916 3398 181944 12310
rect 182008 7342 182036 71726
rect 182836 69086 182864 71726
rect 183480 71726 183525 71754
rect 184194 71754 184222 72012
rect 184892 71754 184920 72012
rect 184194 71726 184244 71754
rect 182088 69080 182140 69086
rect 182088 69022 182140 69028
rect 182824 69080 182876 69086
rect 182824 69022 182876 69028
rect 183376 69080 183428 69086
rect 183376 69022 183428 69028
rect 181996 7336 182048 7342
rect 181996 7278 182048 7284
rect 182100 7274 182128 69022
rect 183388 7410 183416 69022
rect 183480 7478 183508 71726
rect 184216 69086 184244 71726
rect 184768 71726 184920 71754
rect 185590 71754 185618 72012
rect 186288 71754 186316 72012
rect 186986 71754 187014 72012
rect 185590 71726 185624 71754
rect 186288 71726 186360 71754
rect 184204 69080 184256 69086
rect 184204 69022 184256 69028
rect 183744 9308 183796 9314
rect 183744 9250 183796 9256
rect 183468 7472 183520 7478
rect 183468 7414 183520 7420
rect 183376 7404 183428 7410
rect 183376 7346 183428 7352
rect 182088 7268 182140 7274
rect 182088 7210 182140 7216
rect 182548 4752 182600 4758
rect 182548 4694 182600 4700
rect 181444 3392 181496 3398
rect 181444 3334 181496 3340
rect 181904 3392 181956 3398
rect 181904 3334 181956 3340
rect 181456 480 181484 3334
rect 182560 480 182588 4694
rect 183756 480 183784 9250
rect 184768 8294 184796 71726
rect 185596 69086 185624 71726
rect 186332 69154 186360 71726
rect 186976 71726 187014 71754
rect 187683 71754 187711 72012
rect 188381 71754 188409 72012
rect 187683 71726 187740 71754
rect 186320 69148 186372 69154
rect 186320 69090 186372 69096
rect 186976 69086 187004 71726
rect 187712 69154 187740 71726
rect 188356 71726 188409 71754
rect 189079 71754 189107 72012
rect 189777 71754 189805 72012
rect 190475 71754 190503 72012
rect 189079 71726 189120 71754
rect 189777 71726 189856 71754
rect 187608 69148 187660 69154
rect 187608 69090 187660 69096
rect 187700 69148 187752 69154
rect 187700 69090 187752 69096
rect 184848 69080 184900 69086
rect 184848 69022 184900 69028
rect 185584 69080 185636 69086
rect 185584 69022 185636 69028
rect 186228 69080 186280 69086
rect 186228 69022 186280 69028
rect 186964 69080 187016 69086
rect 186964 69022 187016 69028
rect 187516 69080 187568 69086
rect 187516 69022 187568 69028
rect 184756 8288 184808 8294
rect 184756 8230 184808 8236
rect 184860 7546 184888 69022
rect 186240 8226 186268 69022
rect 187332 10804 187384 10810
rect 187332 10746 187384 10752
rect 186228 8220 186280 8226
rect 186228 8162 186280 8168
rect 184848 7540 184900 7546
rect 184848 7482 184900 7488
rect 186136 5500 186188 5506
rect 186136 5442 186188 5448
rect 184940 3868 184992 3874
rect 184940 3810 184992 3816
rect 184952 480 184980 3810
rect 186148 480 186176 5442
rect 187344 480 187372 10746
rect 187528 8090 187556 69022
rect 187620 8158 187648 69090
rect 188356 69086 188384 71726
rect 189092 69154 189120 71726
rect 188896 69148 188948 69154
rect 188896 69090 188948 69096
rect 189080 69148 189132 69154
rect 189080 69090 189132 69096
rect 188344 69080 188396 69086
rect 188344 69022 188396 69028
rect 187608 8152 187660 8158
rect 187608 8094 187660 8100
rect 187516 8084 187568 8090
rect 187516 8026 187568 8032
rect 188908 8022 188936 69090
rect 189828 69086 189856 71726
rect 190472 71726 190503 71754
rect 191172 71754 191200 72012
rect 191870 71754 191898 72012
rect 191172 71726 191236 71754
rect 190472 69154 190500 71726
rect 190276 69148 190328 69154
rect 190276 69090 190328 69096
rect 190460 69148 190512 69154
rect 190460 69090 190512 69096
rect 188988 69080 189040 69086
rect 188988 69022 189040 69028
rect 189816 69080 189868 69086
rect 189816 69022 189868 69028
rect 188896 8016 188948 8022
rect 188896 7958 188948 7964
rect 189000 7954 189028 69022
rect 188988 7948 189040 7954
rect 188988 7890 189040 7896
rect 190288 7886 190316 69090
rect 191208 69086 191236 71726
rect 191852 71726 191898 71754
rect 192568 71754 192596 72012
rect 193266 71754 193294 72012
rect 193964 71754 193992 72012
rect 194661 71754 194689 72012
rect 195359 71754 195387 72012
rect 192568 71726 192616 71754
rect 193266 71726 193352 71754
rect 193964 71726 193996 71754
rect 194661 71726 194732 71754
rect 191656 69148 191708 69154
rect 191656 69090 191708 69096
rect 190368 69080 190420 69086
rect 190368 69022 190420 69028
rect 191196 69080 191248 69086
rect 191196 69022 191248 69028
rect 190276 7880 190328 7886
rect 190276 7822 190328 7828
rect 190380 7818 190408 69022
rect 191564 10872 191616 10878
rect 191564 10814 191616 10820
rect 190368 7812 190420 7818
rect 190368 7754 190420 7760
rect 189724 5432 189776 5438
rect 189724 5374 189776 5380
rect 188528 4004 188580 4010
rect 188528 3946 188580 3952
rect 188540 480 188568 3946
rect 189736 480 189764 5374
rect 191576 3398 191604 10814
rect 191668 7750 191696 69090
rect 191852 69086 191880 71726
rect 191748 69080 191800 69086
rect 191748 69022 191800 69028
rect 191840 69080 191892 69086
rect 191840 69022 191892 69028
rect 191656 7744 191708 7750
rect 191656 7686 191708 7692
rect 191760 7682 191788 69022
rect 192588 67046 192616 71726
rect 193324 69698 193352 71726
rect 193312 69692 193364 69698
rect 193312 69634 193364 69640
rect 193128 69080 193180 69086
rect 193128 69022 193180 69028
rect 192576 67040 192628 67046
rect 192576 66982 192628 66988
rect 191748 7676 191800 7682
rect 191748 7618 191800 7624
rect 193140 7614 193168 69022
rect 193968 68474 193996 71726
rect 194704 69154 194732 71726
rect 195348 71726 195387 71754
rect 196057 71754 196085 72012
rect 196755 71754 196783 72012
rect 196057 71726 196112 71754
rect 194692 69148 194744 69154
rect 194692 69090 194744 69096
rect 195348 69086 195376 71726
rect 196084 69154 196112 71726
rect 196728 71726 196783 71754
rect 197453 71754 197481 72012
rect 198150 71754 198178 72012
rect 198848 71754 198876 72012
rect 197453 71726 197492 71754
rect 198150 71726 198228 71754
rect 195888 69148 195940 69154
rect 195888 69090 195940 69096
rect 196072 69148 196124 69154
rect 196072 69090 196124 69096
rect 195336 69080 195388 69086
rect 195336 69022 195388 69028
rect 195796 69080 195848 69086
rect 195796 69022 195848 69028
rect 193956 68468 194008 68474
rect 193956 68410 194008 68416
rect 195244 17400 195296 17406
rect 195244 17342 195296 17348
rect 193128 7608 193180 7614
rect 193128 7550 193180 7556
rect 193220 5364 193272 5370
rect 193220 5306 193272 5312
rect 192024 3936 192076 3942
rect 192024 3878 192076 3884
rect 190828 3392 190880 3398
rect 190828 3334 190880 3340
rect 191564 3392 191616 3398
rect 191564 3334 191616 3340
rect 190840 480 190868 3334
rect 192036 480 192064 3878
rect 193232 480 193260 5306
rect 194416 4208 194468 4214
rect 194416 4150 194468 4156
rect 194428 480 194456 4150
rect 195256 4010 195284 17342
rect 195336 14816 195388 14822
rect 195336 14758 195388 14764
rect 195244 4004 195296 4010
rect 195244 3946 195296 3952
rect 195348 3806 195376 14758
rect 195808 14482 195836 69022
rect 195796 14476 195848 14482
rect 195796 14418 195848 14424
rect 195612 13660 195664 13666
rect 195612 13602 195664 13608
rect 195336 3800 195388 3806
rect 195336 3742 195388 3748
rect 195624 480 195652 13602
rect 195900 13258 195928 69090
rect 196728 69086 196756 71726
rect 197176 69148 197228 69154
rect 197176 69090 197228 69096
rect 196716 69080 196768 69086
rect 196716 69022 196768 69028
rect 196624 16176 196676 16182
rect 196624 16118 196676 16124
rect 195888 13252 195940 13258
rect 195888 13194 195940 13200
rect 196636 3874 196664 16118
rect 197188 15910 197216 69090
rect 197268 69080 197320 69086
rect 197268 69022 197320 69028
rect 197176 15904 197228 15910
rect 197176 15846 197228 15852
rect 197280 11830 197308 69022
rect 197464 65618 197492 71726
rect 198004 69216 198056 69222
rect 198004 69158 198056 69164
rect 197452 65612 197504 65618
rect 197452 65554 197504 65560
rect 197268 11824 197320 11830
rect 197268 11766 197320 11772
rect 196808 5296 196860 5302
rect 196808 5238 196860 5244
rect 196624 3868 196676 3874
rect 196624 3810 196676 3816
rect 196820 480 196848 5238
rect 198016 4214 198044 69158
rect 198200 69086 198228 71726
rect 198844 71726 198876 71754
rect 199546 71754 199574 72012
rect 200244 71754 200272 72012
rect 199546 71726 199608 71754
rect 198844 69154 198872 71726
rect 198832 69148 198884 69154
rect 198832 69090 198884 69096
rect 199580 69086 199608 71726
rect 200224 71726 200272 71754
rect 200942 71754 200970 72012
rect 201639 71754 201667 72012
rect 202337 71754 202365 72012
rect 203035 71754 203063 72012
rect 203733 71754 203761 72012
rect 200942 71726 201356 71754
rect 201639 71726 201724 71754
rect 202337 71726 202736 71754
rect 203035 71726 203104 71754
rect 199936 69148 199988 69154
rect 199936 69090 199988 69096
rect 198188 69080 198240 69086
rect 198188 69022 198240 69028
rect 198648 69080 198700 69086
rect 198648 69022 198700 69028
rect 199568 69080 199620 69086
rect 199568 69022 199620 69028
rect 198556 18828 198608 18834
rect 198556 18770 198608 18776
rect 198004 4208 198056 4214
rect 198004 4150 198056 4156
rect 198568 3398 198596 18770
rect 198660 13190 198688 69022
rect 198648 13184 198700 13190
rect 198648 13126 198700 13132
rect 199948 9586 199976 69090
rect 200224 69086 200252 71726
rect 200028 69080 200080 69086
rect 200028 69022 200080 69028
rect 200212 69080 200264 69086
rect 200212 69022 200264 69028
rect 199936 9580 199988 9586
rect 199936 9522 199988 9528
rect 200040 9450 200068 69022
rect 200028 9444 200080 9450
rect 200028 9386 200080 9392
rect 201328 9178 201356 71726
rect 201696 69086 201724 71726
rect 201408 69080 201460 69086
rect 201408 69022 201460 69028
rect 201684 69080 201736 69086
rect 201684 69022 201736 69028
rect 201420 9382 201448 69022
rect 202604 18692 202656 18698
rect 202604 18634 202656 18640
rect 202512 10940 202564 10946
rect 202512 10882 202564 10888
rect 201408 9376 201460 9382
rect 201408 9318 201460 9324
rect 201316 9172 201368 9178
rect 201316 9114 201368 9120
rect 200304 5228 200356 5234
rect 200304 5170 200356 5176
rect 199108 3800 199160 3806
rect 199108 3742 199160 3748
rect 197912 3392 197964 3398
rect 197912 3334 197964 3340
rect 198556 3392 198608 3398
rect 198556 3334 198608 3340
rect 197924 480 197952 3334
rect 199120 480 199148 3742
rect 200316 480 200344 5170
rect 202524 3398 202552 10882
rect 202616 6914 202644 18634
rect 202708 9042 202736 71726
rect 203076 69086 203104 71726
rect 203720 71726 203761 71754
rect 204431 71754 204459 72012
rect 205128 71754 205156 72012
rect 204431 71726 204484 71754
rect 203720 69154 203748 71726
rect 203708 69148 203760 69154
rect 203708 69090 203760 69096
rect 202788 69080 202840 69086
rect 202788 69022 202840 69028
rect 203064 69080 203116 69086
rect 203064 69022 203116 69028
rect 204168 69080 204220 69086
rect 204168 69022 204220 69028
rect 202800 9110 202828 69022
rect 202788 9104 202840 9110
rect 202788 9046 202840 9052
rect 202696 9036 202748 9042
rect 202696 8978 202748 8984
rect 204180 8974 204208 69022
rect 204456 68406 204484 71726
rect 205100 71726 205156 71754
rect 205826 71754 205854 72012
rect 206524 71754 206552 72012
rect 207222 71754 207250 72012
rect 205826 71726 205864 71754
rect 206524 71726 206968 71754
rect 204904 69760 204956 69766
rect 204956 69708 205036 69714
rect 204904 69702 205036 69708
rect 204916 69686 205036 69702
rect 205100 69698 205128 71726
rect 204904 69352 204956 69358
rect 204904 69294 204956 69300
rect 204444 68400 204496 68406
rect 204444 68342 204496 68348
rect 204168 8968 204220 8974
rect 204168 8910 204220 8916
rect 202616 6886 202736 6914
rect 201500 3392 201552 3398
rect 201500 3334 201552 3340
rect 202512 3392 202564 3398
rect 202512 3334 202564 3340
rect 201512 480 201540 3334
rect 202708 480 202736 6886
rect 204916 6730 204944 69294
rect 204904 6724 204956 6730
rect 204904 6666 204956 6672
rect 205008 6118 205036 69686
rect 205088 69692 205140 69698
rect 205088 69634 205140 69640
rect 205836 66978 205864 71726
rect 206284 69420 206336 69426
rect 206284 69362 206336 69368
rect 205824 66972 205876 66978
rect 205824 66914 205876 66920
rect 206296 6866 206324 69362
rect 206376 14884 206428 14890
rect 206376 14826 206428 14832
rect 206284 6860 206336 6866
rect 206284 6802 206336 6808
rect 205088 6792 205140 6798
rect 205088 6734 205140 6740
rect 204996 6112 205048 6118
rect 204996 6054 205048 6060
rect 203892 5160 203944 5166
rect 203892 5102 203944 5108
rect 203904 480 203932 5102
rect 205100 480 205128 6734
rect 206388 3942 206416 14826
rect 206940 13122 206968 71726
rect 207216 71726 207250 71754
rect 207920 71754 207948 72012
rect 208617 71754 208645 72012
rect 207920 71726 207980 71754
rect 207216 69358 207244 71726
rect 207204 69352 207256 69358
rect 207204 69294 207256 69300
rect 207952 69154 207980 71726
rect 208596 71726 208645 71754
rect 209315 71754 209343 72012
rect 210013 71754 210041 72012
rect 210711 71754 210739 72012
rect 211409 71754 211437 72012
rect 212106 71754 212134 72012
rect 212804 71754 212832 72012
rect 213502 71754 213530 72012
rect 214200 71754 214228 72012
rect 214898 71754 214926 72012
rect 215595 71754 215623 72012
rect 209315 71726 209360 71754
rect 210013 71726 210096 71754
rect 210711 71726 211108 71754
rect 211409 71726 211476 71754
rect 212106 71726 212488 71754
rect 212804 71726 212856 71754
rect 213502 71726 213776 71754
rect 214200 71726 214236 71754
rect 214898 71726 215248 71754
rect 208596 69766 208624 71726
rect 208584 69760 208636 69766
rect 208584 69702 208636 69708
rect 209136 69284 209188 69290
rect 209136 69226 209188 69232
rect 207940 69148 207992 69154
rect 207940 69090 207992 69096
rect 209044 67244 209096 67250
rect 209044 67186 209096 67192
rect 206928 13116 206980 13122
rect 206928 13058 206980 13064
rect 207388 5092 207440 5098
rect 207388 5034 207440 5040
rect 206376 3936 206428 3942
rect 206376 3878 206428 3884
rect 206192 3868 206244 3874
rect 206192 3810 206244 3816
rect 206204 480 206232 3810
rect 207400 480 207428 5034
rect 209056 3806 209084 67186
rect 209148 10742 209176 69226
rect 209332 66910 209360 71726
rect 209688 69420 209740 69426
rect 209688 69362 209740 69368
rect 209320 66904 209372 66910
rect 209320 66846 209372 66852
rect 209136 10736 209188 10742
rect 209136 10678 209188 10684
rect 209044 3800 209096 3806
rect 209044 3742 209096 3748
rect 209700 3398 209728 69362
rect 210068 69086 210096 71726
rect 210056 69080 210108 69086
rect 210056 69022 210108 69028
rect 210976 69080 211028 69086
rect 210976 69022 211028 69028
rect 210988 6914 211016 69022
rect 210896 6886 211016 6914
rect 210896 4350 210924 6886
rect 210976 5024 211028 5030
rect 210976 4966 211028 4972
rect 210884 4344 210936 4350
rect 210884 4286 210936 4292
rect 209780 3936 209832 3942
rect 209780 3878 209832 3884
rect 208584 3392 208636 3398
rect 208584 3334 208636 3340
rect 209688 3392 209740 3398
rect 209688 3334 209740 3340
rect 208596 480 208624 3334
rect 209792 480 209820 3878
rect 210988 480 211016 4966
rect 211080 4418 211108 71726
rect 211448 69086 211476 71726
rect 211436 69080 211488 69086
rect 211436 69022 211488 69028
rect 212356 69080 212408 69086
rect 212356 69022 212408 69028
rect 212172 5908 212224 5914
rect 212172 5850 212224 5856
rect 211068 4412 211120 4418
rect 211068 4354 211120 4360
rect 212184 480 212212 5850
rect 212368 4486 212396 69022
rect 212460 4554 212488 71726
rect 212828 69086 212856 71726
rect 213644 69148 213696 69154
rect 213644 69090 213696 69096
rect 212816 69080 212868 69086
rect 212816 69022 212868 69028
rect 213656 68338 213684 69090
rect 213644 68332 213696 68338
rect 213644 68274 213696 68280
rect 213748 4690 213776 71726
rect 214208 69086 214236 71726
rect 213828 69080 213880 69086
rect 213828 69022 213880 69028
rect 214196 69080 214248 69086
rect 214196 69022 214248 69028
rect 215116 69080 215168 69086
rect 215116 69022 215168 69028
rect 213736 4684 213788 4690
rect 213736 4626 213788 4632
rect 213840 4622 213868 69022
rect 214472 4956 214524 4962
rect 214472 4898 214524 4904
rect 213828 4616 213880 4622
rect 213828 4558 213880 4564
rect 212448 4548 212500 4554
rect 212448 4490 212500 4496
rect 212356 4480 212408 4486
rect 212356 4422 212408 4428
rect 213368 3800 213420 3806
rect 213368 3742 213420 3748
rect 213380 480 213408 3742
rect 214484 480 214512 4898
rect 215128 4758 215156 69022
rect 215220 5506 215248 71726
rect 215588 71726 215623 71754
rect 216293 71754 216321 72012
rect 216991 71754 217019 72012
rect 216293 71726 216628 71754
rect 215588 69086 215616 71726
rect 215576 69080 215628 69086
rect 215576 69022 215628 69028
rect 216496 69080 216548 69086
rect 216496 69022 216548 69028
rect 215668 9648 215720 9654
rect 215668 9590 215720 9596
rect 215208 5500 215260 5506
rect 215208 5442 215260 5448
rect 215116 4752 215168 4758
rect 215116 4694 215168 4700
rect 215680 480 215708 9590
rect 216508 5438 216536 69022
rect 216496 5432 216548 5438
rect 216496 5374 216548 5380
rect 216600 5370 216628 71726
rect 216968 71726 217019 71754
rect 217689 71754 217717 72012
rect 218387 71754 218415 72012
rect 217689 71726 218008 71754
rect 218387 71726 218468 71754
rect 216968 69086 216996 71726
rect 216956 69080 217008 69086
rect 216956 69022 217008 69028
rect 217876 69080 217928 69086
rect 217876 69022 217928 69028
rect 216588 5364 216640 5370
rect 216588 5306 216640 5312
rect 217888 5302 217916 69022
rect 217876 5296 217928 5302
rect 217876 5238 217928 5244
rect 217980 5234 218008 71726
rect 218440 69086 218468 71726
rect 218428 69080 218480 69086
rect 218428 69022 218480 69028
rect 218980 69080 219032 69086
rect 218980 69022 219032 69028
rect 218992 64874 219020 69022
rect 219084 68490 219112 72012
rect 219782 71754 219810 72012
rect 220480 71754 220508 72012
rect 221178 71754 221206 72012
rect 221876 71754 221904 72012
rect 222573 71890 222601 72012
rect 222573 71862 222608 71890
rect 219782 71726 219848 71754
rect 220480 71726 220768 71754
rect 221178 71726 221228 71754
rect 221876 71726 222056 71754
rect 219820 69086 219848 71726
rect 219808 69080 219860 69086
rect 219808 69022 219860 69028
rect 220636 69080 220688 69086
rect 220636 69022 220688 69028
rect 219084 68462 219388 68490
rect 218992 64846 219296 64874
rect 219268 6914 219296 64846
rect 219176 6886 219296 6914
rect 217968 5228 218020 5234
rect 217968 5170 218020 5176
rect 219176 5166 219204 6886
rect 219256 5976 219308 5982
rect 219256 5918 219308 5924
rect 219164 5160 219216 5166
rect 219164 5102 219216 5108
rect 218060 4888 218112 4894
rect 218060 4830 218112 4836
rect 216864 4072 216916 4078
rect 216864 4014 216916 4020
rect 216876 480 216904 4014
rect 218072 480 218100 4830
rect 219268 480 219296 5918
rect 219360 5098 219388 68462
rect 219348 5092 219400 5098
rect 219348 5034 219400 5040
rect 220648 5030 220676 69022
rect 220636 5024 220688 5030
rect 220636 4966 220688 4972
rect 220740 4962 220768 71726
rect 221200 69086 221228 71726
rect 221188 69080 221240 69086
rect 221188 69022 221240 69028
rect 220728 4956 220780 4962
rect 220728 4898 220780 4904
rect 222028 4826 222056 71726
rect 222108 69080 222160 69086
rect 222108 69022 222160 69028
rect 222120 4894 222148 69022
rect 222580 65550 222608 71862
rect 223271 71754 223299 72012
rect 223969 71754 223997 72012
rect 222764 71726 223299 71754
rect 223960 71726 223997 71754
rect 224667 71754 224695 72012
rect 225365 71754 225393 72012
rect 224667 71726 224724 71754
rect 222568 65544 222620 65550
rect 222568 65486 222620 65492
rect 222764 64874 222792 71726
rect 223960 69834 223988 71726
rect 224696 70038 224724 71726
rect 225340 71726 225393 71754
rect 226062 71754 226090 72012
rect 226760 71754 226788 72012
rect 227458 71754 227486 72012
rect 228156 71754 228184 72012
rect 228854 71754 228882 72012
rect 226062 71726 226104 71754
rect 225340 70174 225368 71726
rect 226076 70310 226104 71726
rect 226720 71726 226788 71754
rect 227456 71726 227486 71754
rect 227824 71726 228184 71754
rect 228836 71726 228882 71754
rect 229551 71754 229579 72012
rect 230249 71754 230277 72012
rect 229551 71726 229600 71754
rect 226064 70304 226116 70310
rect 226064 70246 226116 70252
rect 226720 70242 226748 71726
rect 227456 70378 227484 71726
rect 227444 70372 227496 70378
rect 227444 70314 227496 70320
rect 226708 70236 226760 70242
rect 226708 70178 226760 70184
rect 225328 70168 225380 70174
rect 225328 70110 225380 70116
rect 224684 70032 224736 70038
rect 224684 69974 224736 69980
rect 223948 69828 224000 69834
rect 223948 69770 224000 69776
rect 227628 69624 227680 69630
rect 227628 69566 227680 69572
rect 224224 69556 224276 69562
rect 224224 69498 224276 69504
rect 222844 69284 222896 69290
rect 222844 69226 222896 69232
rect 222212 64846 222792 64874
rect 222212 9246 222240 64846
rect 222856 9518 222884 69226
rect 222936 18760 222988 18766
rect 222936 18702 222988 18708
rect 222844 9512 222896 9518
rect 222844 9454 222896 9460
rect 222200 9240 222252 9246
rect 222200 9182 222252 9188
rect 222752 9240 222804 9246
rect 222752 9182 222804 9188
rect 222108 4888 222160 4894
rect 222108 4830 222160 4836
rect 221556 4820 221608 4826
rect 221556 4762 221608 4768
rect 222016 4820 222068 4826
rect 222016 4762 222068 4768
rect 220452 2916 220504 2922
rect 220452 2858 220504 2864
rect 220464 480 220492 2858
rect 221568 480 221596 4762
rect 222764 480 222792 9182
rect 222948 2922 222976 18702
rect 224236 6050 224264 69498
rect 226984 69488 227036 69494
rect 226984 69430 227036 69436
rect 224316 69352 224368 69358
rect 224316 69294 224368 69300
rect 224328 11762 224356 69294
rect 224408 16244 224460 16250
rect 224408 16186 224460 16192
rect 224316 11756 224368 11762
rect 224316 11698 224368 11704
rect 224224 6044 224276 6050
rect 224224 5986 224276 5992
rect 223948 4004 224000 4010
rect 223948 3946 224000 3952
rect 222936 2916 222988 2922
rect 222936 2858 222988 2864
rect 223960 480 223988 3946
rect 224420 3874 224448 16186
rect 226996 11694 227024 69430
rect 227076 22772 227128 22778
rect 227076 22714 227128 22720
rect 226984 11688 227036 11694
rect 226984 11630 227036 11636
rect 225144 4276 225196 4282
rect 225144 4218 225196 4224
rect 224408 3868 224460 3874
rect 224408 3810 224460 3816
rect 225156 480 225184 4218
rect 227088 4078 227116 22714
rect 227076 4072 227128 4078
rect 227076 4014 227128 4020
rect 227536 3936 227588 3942
rect 227536 3878 227588 3884
rect 226340 3392 226392 3398
rect 226340 3334 226392 3340
rect 226352 480 226380 3334
rect 227548 480 227576 3878
rect 227640 3398 227668 69566
rect 227824 12102 227852 71726
rect 228364 69828 228416 69834
rect 228364 69770 228416 69776
rect 227812 12096 227864 12102
rect 227812 12038 227864 12044
rect 228376 10674 228404 69770
rect 228836 69562 228864 71726
rect 228824 69556 228876 69562
rect 228824 69498 228876 69504
rect 229572 68542 229600 71726
rect 230216 71726 230277 71754
rect 230480 71800 230532 71806
rect 230947 71754 230975 72012
rect 231645 71806 231673 72012
rect 230480 71742 230532 71748
rect 230216 69834 230244 71726
rect 230204 69828 230256 69834
rect 230204 69770 230256 69776
rect 229560 68536 229612 68542
rect 229560 68478 229612 68484
rect 228456 44872 228508 44878
rect 228456 44814 228508 44820
rect 228364 10668 228416 10674
rect 228364 10610 228416 10616
rect 228468 3874 228496 44814
rect 230492 12170 230520 71742
rect 230584 71726 230975 71754
rect 231633 71800 231685 71806
rect 232343 71754 232371 72012
rect 233040 71754 233068 72012
rect 233738 71890 233766 72012
rect 231633 71742 231685 71748
rect 231872 71726 232371 71754
rect 232424 71726 233068 71754
rect 233252 71862 233766 71890
rect 230584 14550 230612 71726
rect 231124 70168 231176 70174
rect 231124 70110 231176 70116
rect 230572 14544 230624 14550
rect 230572 14486 230624 14492
rect 230480 12164 230532 12170
rect 230480 12106 230532 12112
rect 228732 6112 228784 6118
rect 228732 6054 228784 6060
rect 229836 6112 229888 6118
rect 229836 6054 229888 6060
rect 228456 3868 228508 3874
rect 228456 3810 228508 3816
rect 227628 3392 227680 3398
rect 227628 3334 227680 3340
rect 228744 480 228772 6054
rect 229848 480 229876 6054
rect 231136 5914 231164 70110
rect 231216 14952 231268 14958
rect 231216 14894 231268 14900
rect 231124 5908 231176 5914
rect 231124 5850 231176 5856
rect 231228 3942 231256 14894
rect 231872 13734 231900 71726
rect 232424 64874 232452 71726
rect 233252 69290 233280 71862
rect 234436 71754 234464 72012
rect 233344 71726 234464 71754
rect 234712 71800 234764 71806
rect 235134 71754 235162 72012
rect 235832 71806 235860 72012
rect 234712 71742 234764 71748
rect 233240 69284 233292 69290
rect 233240 69226 233292 69232
rect 232504 69080 232556 69086
rect 232504 69022 232556 69028
rect 231964 64846 232452 64874
rect 231964 17474 231992 64846
rect 231952 17468 232004 17474
rect 231952 17410 232004 17416
rect 231860 13728 231912 13734
rect 231860 13670 231912 13676
rect 231768 13592 231820 13598
rect 231768 13534 231820 13540
rect 231216 3936 231268 3942
rect 231216 3878 231268 3884
rect 231780 3398 231808 13534
rect 232516 10810 232544 69022
rect 232596 17468 232648 17474
rect 232596 17410 232648 17416
rect 232504 10804 232556 10810
rect 232504 10746 232556 10752
rect 232228 6860 232280 6866
rect 232228 6802 232280 6808
rect 231032 3392 231084 3398
rect 231032 3334 231084 3340
rect 231768 3392 231820 3398
rect 231768 3334 231820 3340
rect 231044 480 231072 3334
rect 232240 480 232268 6802
rect 232608 3806 232636 17410
rect 233344 9314 233372 71726
rect 234528 70032 234580 70038
rect 234528 69974 234580 69980
rect 233332 9308 233384 9314
rect 233332 9250 233384 9256
rect 232596 3800 232648 3806
rect 232596 3742 232648 3748
rect 234540 3398 234568 69974
rect 234724 10878 234752 71742
rect 235092 71726 235162 71754
rect 235820 71800 235872 71806
rect 235820 71742 235872 71748
rect 236092 71800 236144 71806
rect 236529 71754 236557 72012
rect 237227 71806 237255 72012
rect 236092 71742 236144 71748
rect 235092 69086 235120 71726
rect 235080 69080 235132 69086
rect 235080 69022 235132 69028
rect 235908 50380 235960 50386
rect 235908 50322 235960 50328
rect 234712 10872 234764 10878
rect 234712 10814 234764 10820
rect 235816 6656 235868 6662
rect 235816 6598 235868 6604
rect 233424 3392 233476 3398
rect 233424 3334 233476 3340
rect 234528 3392 234580 3398
rect 234528 3334 234580 3340
rect 234620 3392 234672 3398
rect 234620 3334 234672 3340
rect 233436 480 233464 3334
rect 234632 480 234660 3334
rect 235828 480 235856 6598
rect 235920 3398 235948 50322
rect 236104 18834 236132 71742
rect 236472 71726 236557 71754
rect 237215 71800 237267 71806
rect 237215 71742 237267 71748
rect 237380 71800 237432 71806
rect 237925 71754 237953 72012
rect 238623 71806 238651 72012
rect 237380 71742 237432 71748
rect 236472 69222 236500 71726
rect 236460 69216 236512 69222
rect 236460 69158 236512 69164
rect 236092 18828 236144 18834
rect 236092 18770 236144 18776
rect 237392 6798 237420 71742
rect 237484 71726 237953 71754
rect 238611 71800 238663 71806
rect 238611 71742 238663 71748
rect 239321 71754 239349 72012
rect 240018 71754 240046 72012
rect 239321 71726 239352 71754
rect 237484 10946 237512 71726
rect 239324 69426 239352 71726
rect 239968 71726 240046 71754
rect 240140 71800 240192 71806
rect 240716 71754 240744 72012
rect 241414 71806 241442 72012
rect 240140 71742 240192 71748
rect 239968 70174 239996 71726
rect 239956 70168 240008 70174
rect 239956 70110 240008 70116
rect 239312 69420 239364 69426
rect 239312 69362 239364 69368
rect 238024 25560 238076 25566
rect 238024 25502 238076 25508
rect 237472 10940 237524 10946
rect 237472 10882 237524 10888
rect 237380 6792 237432 6798
rect 237380 6734 237432 6740
rect 237012 6656 237064 6662
rect 237012 6598 237064 6604
rect 235908 3392 235960 3398
rect 235908 3334 235960 3340
rect 237024 480 237052 6598
rect 238036 4010 238064 25502
rect 239312 6724 239364 6730
rect 239312 6666 239364 6672
rect 238024 4004 238076 4010
rect 238024 3946 238076 3952
rect 238116 3800 238168 3806
rect 238116 3742 238168 3748
rect 238128 480 238156 3742
rect 239324 480 239352 6666
rect 240152 5982 240180 71742
rect 240244 71726 240744 71754
rect 241402 71800 241454 71806
rect 242112 71754 242140 72012
rect 241402 71742 241454 71748
rect 241624 71726 242140 71754
rect 242810 71754 242838 72012
rect 243507 71754 243535 72012
rect 244205 71754 244233 72012
rect 244903 71754 244931 72012
rect 245601 71754 245629 72012
rect 246299 71754 246327 72012
rect 246996 71754 247024 72012
rect 242810 71726 242848 71754
rect 240244 9654 240272 71726
rect 240232 9648 240284 9654
rect 240232 9590 240284 9596
rect 240508 9648 240560 9654
rect 240508 9590 240560 9596
rect 240140 5976 240192 5982
rect 240140 5918 240192 5924
rect 240520 480 240548 9590
rect 241624 9246 241652 71726
rect 242820 69834 242848 71726
rect 243464 71726 243535 71754
rect 244200 71726 244233 71754
rect 244292 71726 244931 71754
rect 245580 71726 245629 71754
rect 245672 71726 246327 71754
rect 246960 71726 247024 71754
rect 247694 71754 247722 72012
rect 248392 71754 248420 72012
rect 249090 71754 249118 72012
rect 247694 71726 247724 71754
rect 248392 71726 248460 71754
rect 242808 69828 242860 69834
rect 242808 69770 242860 69776
rect 243464 69086 243492 71726
rect 244200 70038 244228 71726
rect 244188 70032 244240 70038
rect 244188 69974 244240 69980
rect 242164 69080 242216 69086
rect 242164 69022 242216 69028
rect 243452 69080 243504 69086
rect 243452 69022 243504 69028
rect 241612 9240 241664 9246
rect 241612 9182 241664 9188
rect 242176 6118 242204 69022
rect 242256 17604 242308 17610
rect 242256 17546 242308 17552
rect 242164 6112 242216 6118
rect 242164 6054 242216 6060
rect 242268 3806 242296 17546
rect 244292 6662 244320 71726
rect 245580 68542 245608 71726
rect 244372 68536 244424 68542
rect 244372 68478 244424 68484
rect 245568 68536 245620 68542
rect 245568 68478 245620 68484
rect 244384 9654 244412 68478
rect 244372 9648 244424 9654
rect 244372 9590 244424 9596
rect 244280 6656 244332 6662
rect 244280 6598 244332 6604
rect 242900 6588 242952 6594
rect 242900 6530 242952 6536
rect 242256 3800 242308 3806
rect 242256 3742 242308 3748
rect 241702 3632 241758 3641
rect 241702 3567 241758 3576
rect 241716 480 241744 3567
rect 242912 480 242940 6530
rect 245672 5574 245700 71726
rect 246396 6044 246448 6050
rect 246396 5986 246448 5992
rect 244096 5568 244148 5574
rect 244096 5510 244148 5516
rect 245660 5568 245712 5574
rect 245660 5510 245712 5516
rect 244108 480 244136 5510
rect 245198 3768 245254 3777
rect 245198 3703 245254 3712
rect 245212 480 245240 3703
rect 246408 480 246436 5986
rect 246960 5574 246988 71726
rect 247696 69630 247724 71726
rect 247684 69624 247736 69630
rect 247684 69566 247736 69572
rect 248432 69154 248460 71726
rect 249076 71726 249118 71754
rect 249788 71754 249816 72012
rect 250485 71754 250513 72012
rect 249788 71726 249840 71754
rect 248972 69624 249024 69630
rect 248972 69566 249024 69572
rect 248420 69148 248472 69154
rect 248420 69090 248472 69096
rect 248984 64874 249012 69566
rect 249076 69086 249104 71726
rect 249708 69148 249760 69154
rect 249708 69090 249760 69096
rect 249064 69080 249116 69086
rect 249064 69022 249116 69028
rect 249616 69080 249668 69086
rect 249616 69022 249668 69028
rect 248984 64846 249104 64874
rect 249076 17950 249104 64846
rect 249064 17944 249116 17950
rect 249064 17886 249116 17892
rect 249628 9246 249656 69022
rect 249616 9240 249668 9246
rect 249616 9182 249668 9188
rect 249720 5574 249748 69090
rect 249812 69086 249840 71726
rect 250456 71726 250513 71754
rect 251183 71754 251211 72012
rect 251881 71754 251909 72012
rect 252579 71754 252607 72012
rect 251183 71726 251220 71754
rect 251881 71726 251956 71754
rect 250352 70168 250404 70174
rect 250352 70110 250404 70116
rect 249800 69080 249852 69086
rect 249800 69022 249852 69028
rect 250364 64874 250392 70110
rect 250456 69834 250484 71726
rect 250444 69828 250496 69834
rect 250444 69770 250496 69776
rect 251192 69154 251220 71726
rect 251180 69148 251232 69154
rect 251180 69090 251232 69096
rect 251928 69086 251956 71726
rect 252572 71726 252607 71754
rect 253277 71754 253305 72012
rect 253974 71754 254002 72012
rect 253277 71726 253336 71754
rect 252572 69154 252600 71726
rect 252468 69148 252520 69154
rect 252468 69090 252520 69096
rect 252560 69148 252612 69154
rect 252560 69090 252612 69096
rect 251088 69080 251140 69086
rect 251088 69022 251140 69028
rect 251916 69080 251968 69086
rect 251916 69022 251968 69028
rect 252376 69080 252428 69086
rect 252376 69022 252428 69028
rect 250364 64846 250484 64874
rect 250456 10606 250484 64846
rect 249984 10600 250036 10606
rect 249984 10542 250036 10548
rect 250444 10600 250496 10606
rect 250444 10542 250496 10548
rect 246948 5568 247000 5574
rect 246948 5510 247000 5516
rect 247592 5568 247644 5574
rect 247592 5510 247644 5516
rect 249708 5568 249760 5574
rect 249708 5510 249760 5516
rect 247604 480 247632 5510
rect 248788 3800 248840 3806
rect 248788 3742 248840 3748
rect 248800 480 248828 3742
rect 249996 480 250024 10542
rect 251100 5914 251128 69022
rect 251180 17944 251232 17950
rect 251180 17886 251232 17892
rect 251088 5908 251140 5914
rect 251088 5850 251140 5856
rect 251192 480 251220 17886
rect 252388 5982 252416 69022
rect 252376 5976 252428 5982
rect 252376 5918 252428 5924
rect 252480 4282 252508 69090
rect 253308 69086 253336 71726
rect 253952 71726 254002 71754
rect 254672 71754 254700 72012
rect 255370 71754 255398 72012
rect 254672 71726 254716 71754
rect 255370 71726 255452 71754
rect 253952 69154 253980 71726
rect 253848 69148 253900 69154
rect 253848 69090 253900 69096
rect 253940 69148 253992 69154
rect 253940 69090 253992 69096
rect 253296 69080 253348 69086
rect 253296 69022 253348 69028
rect 253756 69080 253808 69086
rect 253756 69022 253808 69028
rect 253480 10532 253532 10538
rect 253480 10474 253532 10480
rect 252468 4276 252520 4282
rect 252468 4218 252520 4224
rect 252376 3868 252428 3874
rect 252376 3810 252428 3816
rect 252388 480 252416 3810
rect 253492 480 253520 10474
rect 253768 6118 253796 69022
rect 253756 6112 253808 6118
rect 253756 6054 253808 6060
rect 253860 6050 253888 69090
rect 254688 69086 254716 71726
rect 255424 69154 255452 71726
rect 255228 69148 255280 69154
rect 255228 69090 255280 69096
rect 255412 69148 255464 69154
rect 255412 69090 255464 69096
rect 254676 69080 254728 69086
rect 254676 69022 254728 69028
rect 255136 69080 255188 69086
rect 255136 69022 255188 69028
rect 255148 6798 255176 69022
rect 255240 6866 255268 69090
rect 256068 69086 256096 72012
rect 256766 71754 256794 72012
rect 257463 71754 257491 72012
rect 256766 71726 256832 71754
rect 256804 69154 256832 71726
rect 257448 71726 257491 71754
rect 258161 71754 258189 72012
rect 258859 71754 258887 72012
rect 259557 71754 259585 72012
rect 260255 71754 260283 72012
rect 260952 71754 260980 72012
rect 258161 71726 258212 71754
rect 258859 71726 258948 71754
rect 259557 71726 259592 71754
rect 260255 71726 260696 71754
rect 256608 69148 256660 69154
rect 256608 69090 256660 69096
rect 256792 69148 256844 69154
rect 256792 69090 256844 69096
rect 256056 69080 256108 69086
rect 256056 69022 256108 69028
rect 256516 69080 256568 69086
rect 256516 69022 256568 69028
rect 255228 6860 255280 6866
rect 255228 6802 255280 6808
rect 255136 6792 255188 6798
rect 255136 6734 255188 6740
rect 256528 6662 256556 69022
rect 256620 6730 256648 69090
rect 257448 69086 257476 71726
rect 258184 69154 258212 71726
rect 257896 69148 257948 69154
rect 257896 69090 257948 69096
rect 258172 69148 258224 69154
rect 258172 69090 258224 69096
rect 257436 69080 257488 69086
rect 257436 69022 257488 69028
rect 256608 6724 256660 6730
rect 256608 6666 256660 6672
rect 256516 6656 256568 6662
rect 256516 6598 256568 6604
rect 257908 6594 257936 69090
rect 258920 69086 258948 71726
rect 259276 69148 259328 69154
rect 259276 69090 259328 69096
rect 257988 69080 258040 69086
rect 257988 69022 258040 69028
rect 258908 69080 258960 69086
rect 258908 69022 258960 69028
rect 257896 6588 257948 6594
rect 257896 6530 257948 6536
rect 258000 6526 258028 69022
rect 259288 9518 259316 69090
rect 259564 69086 259592 71726
rect 259368 69080 259420 69086
rect 259368 69022 259420 69028
rect 259552 69080 259604 69086
rect 259552 69022 259604 69028
rect 259276 9512 259328 9518
rect 259276 9454 259328 9460
rect 259380 9314 259408 69022
rect 260668 16574 260696 71726
rect 260944 71726 260980 71754
rect 261650 71754 261678 72012
rect 262348 71754 262376 72012
rect 261650 71726 261708 71754
rect 260944 69154 260972 71726
rect 260932 69148 260984 69154
rect 260932 69090 260984 69096
rect 261680 69086 261708 71726
rect 262324 71726 262376 71754
rect 263046 71754 263074 72012
rect 263744 71754 263772 72012
rect 264441 71754 264469 72012
rect 265139 71754 265167 72012
rect 265837 71754 265865 72012
rect 263046 71726 263088 71754
rect 263744 71726 263824 71754
rect 264441 71726 264836 71754
rect 265139 71726 265204 71754
rect 262324 69154 262352 71726
rect 262036 69148 262088 69154
rect 262036 69090 262088 69096
rect 262312 69148 262364 69154
rect 262312 69090 262364 69096
rect 260748 69080 260800 69086
rect 260748 69022 260800 69028
rect 261668 69080 261720 69086
rect 261668 69022 261720 69028
rect 260576 16546 260696 16574
rect 259368 9308 259420 9314
rect 259368 9250 259420 9256
rect 258264 9240 258316 9246
rect 258264 9182 258316 9188
rect 257068 6520 257120 6526
rect 257068 6462 257120 6468
rect 257988 6520 258040 6526
rect 257988 6462 258040 6468
rect 253848 6044 253900 6050
rect 253848 5986 253900 5992
rect 254676 5568 254728 5574
rect 254676 5510 254728 5516
rect 254688 480 254716 5510
rect 255872 3936 255924 3942
rect 255872 3878 255924 3884
rect 255884 480 255912 3878
rect 257080 480 257108 6462
rect 258276 480 258304 9182
rect 260576 8430 260604 16546
rect 260656 10464 260708 10470
rect 260656 10406 260708 10412
rect 260564 8424 260616 8430
rect 260564 8366 260616 8372
rect 259460 4004 259512 4010
rect 259460 3946 259512 3952
rect 259472 480 259500 3946
rect 260668 480 260696 10406
rect 260760 9246 260788 69022
rect 260748 9240 260800 9246
rect 260748 9182 260800 9188
rect 262048 8498 262076 69090
rect 263060 69086 263088 71726
rect 263416 69148 263468 69154
rect 263416 69090 263468 69096
rect 262128 69080 262180 69086
rect 262128 69022 262180 69028
rect 263048 69080 263100 69086
rect 263048 69022 263100 69028
rect 262140 8566 262168 69022
rect 263428 8634 263456 69090
rect 263796 69086 263824 71726
rect 263508 69080 263560 69086
rect 263508 69022 263560 69028
rect 263784 69080 263836 69086
rect 263784 69022 263836 69028
rect 263520 8702 263548 69022
rect 264152 10396 264204 10402
rect 264152 10338 264204 10344
rect 263508 8696 263560 8702
rect 263508 8638 263560 8644
rect 263416 8628 263468 8634
rect 263416 8570 263468 8576
rect 262128 8560 262180 8566
rect 262128 8502 262180 8508
rect 262036 8492 262088 8498
rect 262036 8434 262088 8440
rect 261760 5908 261812 5914
rect 261760 5850 261812 5856
rect 261772 480 261800 5850
rect 262956 4072 263008 4078
rect 262956 4014 263008 4020
rect 262968 480 262996 4014
rect 264164 480 264192 10338
rect 264808 8838 264836 71726
rect 264980 69828 265032 69834
rect 264980 69770 265032 69776
rect 264888 69080 264940 69086
rect 264888 69022 264940 69028
rect 264796 8832 264848 8838
rect 264796 8774 264848 8780
rect 264900 8770 264928 69022
rect 264888 8764 264940 8770
rect 264888 8706 264940 8712
rect 264992 490 265020 69770
rect 265176 69086 265204 71726
rect 265820 71726 265865 71754
rect 266535 71754 266563 72012
rect 267233 71754 267261 72012
rect 267930 71754 267958 72012
rect 268628 71754 268656 72012
rect 269326 71754 269354 72012
rect 266535 71726 266584 71754
rect 267233 71726 267596 71754
rect 267930 71726 267964 71754
rect 268628 71726 268976 71754
rect 265820 70378 265848 71726
rect 265808 70372 265860 70378
rect 265808 70314 265860 70320
rect 266556 69086 266584 71726
rect 265164 69080 265216 69086
rect 265164 69022 265216 69028
rect 266268 69080 266320 69086
rect 266268 69022 266320 69028
rect 266544 69080 266596 69086
rect 266544 69022 266596 69028
rect 266280 8906 266308 69022
rect 267568 15026 267596 71726
rect 267936 69086 267964 71726
rect 267648 69080 267700 69086
rect 267648 69022 267700 69028
rect 267924 69080 267976 69086
rect 267924 69022 267976 69028
rect 267556 15020 267608 15026
rect 267556 14962 267608 14968
rect 267660 12442 267688 69022
rect 268948 21418 268976 71726
rect 269316 71726 269354 71754
rect 270024 71754 270052 72012
rect 270722 71754 270750 72012
rect 270024 71726 270448 71754
rect 269316 69086 269344 71726
rect 269028 69080 269080 69086
rect 269028 69022 269080 69028
rect 269304 69080 269356 69086
rect 269304 69022 269356 69028
rect 270316 69080 270368 69086
rect 270316 69022 270368 69028
rect 268936 21412 268988 21418
rect 268936 21354 268988 21360
rect 267648 12436 267700 12442
rect 267648 12378 267700 12384
rect 267740 12028 267792 12034
rect 267740 11970 267792 11976
rect 266268 8900 266320 8906
rect 266268 8842 266320 8848
rect 266544 4140 266596 4146
rect 266544 4082 266596 4088
rect 265176 598 265388 626
rect 265176 490 265204 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 598
rect 266556 480 266584 4082
rect 267752 480 267780 11970
rect 269040 4282 269068 69022
rect 270328 16386 270356 69022
rect 270316 16380 270368 16386
rect 270316 16322 270368 16328
rect 270420 13734 270448 71726
rect 270696 71726 270750 71754
rect 271419 71754 271447 72012
rect 272117 71754 272145 72012
rect 272815 71754 272843 72012
rect 273513 71754 273541 72012
rect 274211 71754 274239 72012
rect 274908 71754 274936 72012
rect 275606 71754 275634 72012
rect 276304 71754 276332 72012
rect 277002 71754 277030 72012
rect 277700 71754 277728 72012
rect 271419 71726 271828 71754
rect 272117 71726 272196 71754
rect 272815 71726 273208 71754
rect 273513 71726 273576 71754
rect 274211 71726 274588 71754
rect 274908 71726 274956 71754
rect 275606 71726 275968 71754
rect 276304 71726 276336 71754
rect 277002 71726 277348 71754
rect 270696 69086 270724 71726
rect 270684 69080 270736 69086
rect 270684 69022 270736 69028
rect 271696 69080 271748 69086
rect 271696 69022 271748 69028
rect 271708 17542 271736 69022
rect 271696 17536 271748 17542
rect 271696 17478 271748 17484
rect 271800 16318 271828 71726
rect 272168 69494 272196 71726
rect 272156 69488 272208 69494
rect 272156 69430 272208 69436
rect 271788 16312 271840 16318
rect 271788 16254 271840 16260
rect 270408 13728 270460 13734
rect 270408 13670 270460 13676
rect 270776 10328 270828 10334
rect 270776 10270 270828 10276
rect 268844 4276 268896 4282
rect 268844 4218 268896 4224
rect 269028 4276 269080 4282
rect 269028 4218 269080 4224
rect 268856 480 268884 4218
rect 270040 3392 270092 3398
rect 270040 3334 270092 3340
rect 270052 480 270080 3334
rect 270788 490 270816 10270
rect 273180 9790 273208 71726
rect 273548 69086 273576 71726
rect 274364 69488 274416 69494
rect 274364 69430 274416 69436
rect 273536 69080 273588 69086
rect 273536 69022 273588 69028
rect 274376 67318 274404 69430
rect 274456 69080 274508 69086
rect 274456 69022 274508 69028
rect 274364 67312 274416 67318
rect 274364 67254 274416 67260
rect 274468 9858 274496 69022
rect 274560 9926 274588 71726
rect 274928 69086 274956 71726
rect 274916 69080 274968 69086
rect 274916 69022 274968 69028
rect 275836 69080 275888 69086
rect 275836 69022 275888 69028
rect 274824 10736 274876 10742
rect 274824 10678 274876 10684
rect 274548 9920 274600 9926
rect 274548 9862 274600 9868
rect 274456 9852 274508 9858
rect 274456 9794 274508 9800
rect 273168 9784 273220 9790
rect 273168 9726 273220 9732
rect 272432 5976 272484 5982
rect 272432 5918 272484 5924
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
<<<<<<< HEAD
=======
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 5918
rect 273628 3324 273680 3330
rect 273628 3266 273680 3272
rect 273640 480 273668 3266
rect 274836 480 274864 10678
rect 275848 9994 275876 69022
rect 275940 10062 275968 71726
rect 276308 69086 276336 71726
rect 276296 69080 276348 69086
rect 276296 69022 276348 69028
rect 277216 69080 277268 69086
rect 277216 69022 277268 69028
rect 277228 10130 277256 69022
rect 277320 10198 277348 71726
rect 277688 71726 277728 71754
rect 278397 71754 278425 72012
rect 279095 71754 279123 72012
rect 278397 71726 278728 71754
rect 277688 69086 277716 71726
rect 277676 69080 277728 69086
rect 277676 69022 277728 69028
rect 278596 69080 278648 69086
rect 278596 69022 278648 69028
rect 278320 10600 278372 10606
rect 278320 10542 278372 10548
rect 277308 10192 277360 10198
rect 277308 10134 277360 10140
rect 277216 10124 277268 10130
rect 277216 10066 277268 10072
rect 275928 10056 275980 10062
rect 275928 9998 275980 10004
rect 275836 9988 275888 9994
rect 275836 9930 275888 9936
rect 276020 6044 276072 6050
rect 276020 5986 276072 5992
rect 276032 480 276060 5986
rect 277124 3256 277176 3262
rect 277124 3198 277176 3204
rect 277136 480 277164 3198
rect 278332 480 278360 10542
rect 278608 10266 278636 69022
rect 278700 11014 278728 71726
rect 279068 71726 279123 71754
rect 279793 71754 279821 72012
rect 280491 71754 280519 72012
rect 281189 71754 281217 72012
rect 281886 71754 281914 72012
rect 282584 71754 282612 72012
rect 283282 71754 283310 72012
rect 283980 71754 284008 72012
rect 284678 71754 284706 72012
rect 285375 71754 285403 72012
rect 286073 71754 286101 72012
rect 279793 71726 280108 71754
rect 280491 71726 280568 71754
rect 281189 71726 281304 71754
rect 281886 71726 281948 71754
rect 282584 71726 282868 71754
rect 283282 71726 283328 71754
rect 283980 71726 284156 71754
rect 284678 71726 284708 71754
rect 285375 71726 285628 71754
rect 279068 69086 279096 71726
rect 279056 69080 279108 69086
rect 279056 69022 279108 69028
rect 279976 69080 280028 69086
rect 279976 69022 280028 69028
rect 278688 11008 278740 11014
rect 278688 10950 278740 10956
rect 279988 10946 280016 69022
rect 279976 10940 280028 10946
rect 279976 10882 280028 10888
rect 280080 10878 280108 71726
rect 280540 69086 280568 71726
rect 280528 69080 280580 69086
rect 280528 69022 280580 69028
rect 280068 10872 280120 10878
rect 280068 10814 280120 10820
rect 281276 10742 281304 71726
rect 281448 70168 281500 70174
rect 281448 70110 281500 70116
rect 281356 69080 281408 69086
rect 281356 69022 281408 69028
rect 281368 10810 281396 69022
rect 281356 10804 281408 10810
rect 281356 10746 281408 10752
rect 281264 10736 281316 10742
rect 281264 10678 281316 10684
rect 278596 10260 278648 10266
rect 278596 10202 278648 10208
rect 279516 6112 279568 6118
rect 279516 6054 279568 6060
rect 279528 480 279556 6054
rect 281460 3126 281488 70110
rect 281920 69086 281948 71726
rect 281908 69080 281960 69086
rect 281908 69022 281960 69028
rect 282736 69080 282788 69086
rect 282736 69022 282788 69028
rect 281540 11688 281592 11694
rect 281540 11630 281592 11636
rect 280712 3120 280764 3126
rect 280712 3062 280764 3068
rect 281448 3120 281500 3126
rect 281448 3062 281500 3068
rect 280724 480 280752 3062
rect 281552 490 281580 11630
rect 282748 10674 282776 69022
rect 282736 10668 282788 10674
rect 282736 10610 282788 10616
rect 282840 10606 282868 71726
rect 283300 69086 283328 71726
rect 283288 69080 283340 69086
rect 283288 69022 283340 69028
rect 282828 10600 282880 10606
rect 282828 10542 282880 10548
rect 284128 10470 284156 71726
rect 284680 69086 284708 71726
rect 284208 69080 284260 69086
rect 284208 69022 284260 69028
rect 284668 69080 284720 69086
rect 284668 69022 284720 69028
rect 285496 69080 285548 69086
rect 285496 69022 285548 69028
rect 284220 10538 284248 69022
rect 284944 11892 284996 11898
rect 284944 11834 284996 11840
rect 284208 10532 284260 10538
rect 284208 10474 284260 10480
rect 284116 10464 284168 10470
rect 284116 10406 284168 10412
rect 283104 6860 283156 6866
rect 283104 6802 283156 6808
rect 281736 598 281948 626
rect 281736 490 281764 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 6802
rect 284300 3188 284352 3194
rect 284300 3130 284352 3136
rect 284312 480 284340 3130
rect 284956 490 284984 11834
rect 285508 10402 285536 69022
rect 285496 10396 285548 10402
rect 285496 10338 285548 10344
rect 285600 10334 285628 71726
rect 286060 71726 286101 71754
rect 286771 71754 286799 72012
rect 287469 71754 287497 72012
rect 286771 71726 287008 71754
rect 286060 69086 286088 71726
rect 286048 69080 286100 69086
rect 286048 69022 286100 69028
rect 286876 69080 286928 69086
rect 286876 69022 286928 69028
rect 286888 12170 286916 69022
rect 286876 12164 286928 12170
rect 286876 12106 286928 12112
rect 286980 12102 287008 71726
rect 287440 71726 287497 71754
rect 288167 71754 288195 72012
rect 288864 71754 288892 72012
rect 289562 71754 289590 72012
rect 288167 71726 288296 71754
rect 288864 71726 288940 71754
rect 287440 69086 287468 71726
rect 287704 69828 287756 69834
rect 287704 69770 287756 69776
rect 287428 69080 287480 69086
rect 287428 69022 287480 69028
rect 287716 13666 287744 69770
rect 288268 64190 288296 71726
rect 288912 69086 288940 71726
rect 289556 71726 289590 71754
rect 290260 71754 290288 72012
rect 290958 71754 290986 72012
rect 290260 71726 290320 71754
rect 289084 69488 289136 69494
rect 289084 69430 289136 69436
rect 288348 69080 288400 69086
rect 288348 69022 288400 69028
rect 288900 69080 288952 69086
rect 288900 69022 288952 69028
rect 288256 64184 288308 64190
rect 288256 64126 288308 64132
rect 287704 13660 287756 13666
rect 287704 13602 287756 13608
rect 286968 12096 287020 12102
rect 286968 12038 287020 12044
rect 288360 12034 288388 69022
rect 288348 12028 288400 12034
rect 288348 11970 288400 11976
rect 285588 10328 285640 10334
rect 285588 10270 285640 10276
rect 286600 6792 286652 6798
rect 286600 6734 286652 6740
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 6734
rect 289096 6458 289124 69430
rect 289556 65754 289584 71726
rect 290292 69358 290320 71726
rect 290936 71726 290986 71754
rect 291656 71754 291684 72012
rect 292353 71754 292381 72012
rect 293051 71754 293079 72012
rect 293749 71754 293777 72012
rect 294447 71754 294475 72012
rect 291656 71726 291700 71754
rect 292353 71726 292528 71754
rect 293051 71726 293080 71754
rect 293749 71726 293816 71754
rect 290280 69352 290332 69358
rect 290280 69294 290332 69300
rect 290936 69086 290964 71726
rect 291672 70242 291700 71726
rect 291660 70236 291712 70242
rect 291660 70178 291712 70184
rect 291844 69556 291896 69562
rect 291844 69498 291896 69504
rect 289728 69080 289780 69086
rect 289728 69022 289780 69028
rect 290924 69080 290976 69086
rect 290924 69022 290976 69028
rect 289544 65748 289596 65754
rect 289544 65690 289596 65696
rect 289740 24138 289768 69022
rect 289728 24132 289780 24138
rect 289728 24074 289780 24080
rect 291856 12374 291884 69498
rect 292396 69352 292448 69358
rect 292396 69294 292448 69300
rect 292408 67114 292436 69294
rect 292396 67108 292448 67114
rect 292396 67050 292448 67056
rect 292500 14550 292528 71726
rect 293052 69426 293080 71726
rect 293788 69630 293816 71726
rect 294432 71726 294475 71754
rect 295145 71754 295173 72012
rect 295842 71754 295870 72012
rect 295145 71726 295196 71754
rect 294432 70310 294460 71726
rect 294420 70304 294472 70310
rect 294420 70246 294472 70252
rect 295168 70038 295196 71726
rect 295812 71726 295870 71754
rect 296540 71754 296568 72012
rect 297238 71754 297266 72012
rect 297936 71754 297964 72012
rect 296540 71726 296668 71754
rect 297238 71726 297312 71754
rect 295812 70106 295840 71726
rect 295892 70372 295944 70378
rect 295892 70314 295944 70320
rect 295800 70100 295852 70106
rect 295800 70042 295852 70048
rect 295156 70032 295208 70038
rect 295156 69974 295208 69980
rect 293776 69624 293828 69630
rect 293776 69566 293828 69572
rect 293040 69420 293092 69426
rect 293040 69362 293092 69368
rect 295248 69352 295300 69358
rect 295248 69294 295300 69300
rect 293776 69080 293828 69086
rect 293776 69022 293828 69028
rect 293788 65686 293816 69022
rect 293776 65680 293828 65686
rect 293776 65622 293828 65628
rect 292488 14544 292540 14550
rect 292488 14486 292540 14492
rect 291844 12368 291896 12374
rect 291844 12310 291896 12316
rect 290188 6724 290240 6730
rect 290188 6666 290240 6672
rect 289084 6452 289136 6458
rect 289084 6394 289136 6400
rect 288992 6384 289044 6390
rect 288992 6326 289044 6332
rect 287796 3120 287848 3126
rect 287796 3062 287848 3068
rect 287808 480 287836 3062
rect 289004 480 289032 6326
rect 290200 480 290228 6666
rect 293684 6656 293736 6662
rect 293684 6598 293736 6604
rect 292580 6316 292632 6322
rect 292580 6258 292632 6264
rect 291384 2984 291436 2990
rect 291384 2926 291436 2932
rect 291396 480 291424 2926
rect 292592 480 292620 6258
rect 293696 480 293724 6598
rect 294892 598 295104 626
rect 294892 480 294920 598
rect 295076 490 295104 598
rect 295260 490 295288 69294
rect 295904 64874 295932 70314
rect 295984 70304 296036 70310
rect 295984 70246 296036 70252
rect 295996 68542 296024 70246
rect 295984 68536 296036 68542
rect 295984 68478 296036 68484
rect 295904 64846 296024 64874
rect 295996 19990 296024 64846
rect 295984 19984 296036 19990
rect 295984 19926 296036 19932
rect 296640 11898 296668 71726
rect 297284 69086 297312 71726
rect 297928 71726 297964 71754
rect 298634 71754 298662 72012
rect 299331 71754 299359 72012
rect 298634 71726 298692 71754
rect 297272 69080 297324 69086
rect 297272 69022 297324 69028
rect 296628 11892 296680 11898
rect 296628 11834 296680 11840
rect 297272 6588 297324 6594
rect 297272 6530 297324 6536
rect 296076 6248 296128 6254
rect 296076 6190 296128 6196
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295076 462 295288 490
rect 296088 480 296116 6190
rect 297284 480 297312 6530
rect 297928 5778 297956 71726
rect 298664 69086 298692 71726
rect 299216 71726 299359 71754
rect 300029 71754 300057 72012
rect 300727 71754 300755 72012
rect 301425 71754 301453 72012
rect 302123 71754 302151 72012
rect 302820 71754 302848 72012
rect 303518 71754 303546 72012
rect 300029 71726 300072 71754
rect 300727 71726 300808 71754
rect 298008 69080 298060 69086
rect 298008 69022 298060 69028
rect 298652 69080 298704 69086
rect 298652 69022 298704 69028
rect 297916 5772 297968 5778
rect 297916 5714 297968 5720
rect 298020 5710 298048 69022
rect 299216 5914 299244 71726
rect 299388 70372 299440 70378
rect 299388 70314 299440 70320
rect 299296 69080 299348 69086
rect 299296 69022 299348 69028
rect 299204 5908 299256 5914
rect 299204 5850 299256 5856
rect 299308 5846 299336 69022
rect 299296 5840 299348 5846
rect 299296 5782 299348 5788
rect 298008 5704 298060 5710
rect 298008 5646 298060 5652
rect 299400 2990 299428 70314
rect 300044 69086 300072 71726
rect 300032 69080 300084 69086
rect 300032 69022 300084 69028
rect 300676 69080 300728 69086
rect 300676 69022 300728 69028
rect 300688 16574 300716 69022
rect 300596 16546 300716 16574
rect 299664 6180 299716 6186
rect 299664 6122 299716 6128
rect 298468 2984 298520 2990
rect 298468 2926 298520 2932
rect 299388 2984 299440 2990
rect 299388 2926 299440 2932
rect 298480 480 298508 2926
rect 299676 480 299704 6122
rect 300596 5982 300624 16546
rect 300780 6914 300808 71726
rect 301424 71726 301453 71754
rect 302068 71726 302151 71754
rect 302804 71726 302848 71754
rect 303448 71726 303546 71754
rect 304216 71754 304244 72012
rect 304914 71754 304942 72012
rect 305612 71754 305640 72012
rect 306309 71754 306337 72012
rect 304216 71726 304304 71754
rect 304914 71726 304948 71754
rect 305612 71726 305684 71754
rect 301424 69086 301452 71726
rect 301412 69080 301464 69086
rect 301412 69022 301464 69028
rect 300688 6886 300808 6914
rect 300688 6050 300716 6886
rect 302068 6866 302096 71726
rect 302804 69086 302832 71726
rect 302148 69080 302200 69086
rect 302148 69022 302200 69028
rect 302792 69080 302844 69086
rect 302792 69022 302844 69028
rect 302056 6860 302108 6866
rect 302056 6802 302108 6808
rect 300768 6520 300820 6526
rect 300768 6462 300820 6468
rect 300676 6044 300728 6050
rect 300676 5986 300728 5992
rect 300584 5976 300636 5982
rect 300584 5918 300636 5924
rect 300780 480 300808 6462
rect 302160 6118 302188 69022
rect 303160 12300 303212 12306
rect 303160 12242 303212 12248
rect 302148 6112 302200 6118
rect 302148 6054 302200 6060
rect 301964 2984 302016 2990
rect 301964 2926 302016 2932
rect 301976 480 302004 2926
rect 303172 480 303200 12242
rect 303448 6730 303476 71726
rect 304276 69086 304304 71726
rect 303528 69080 303580 69086
rect 303528 69022 303580 69028
rect 304264 69080 304316 69086
rect 304264 69022 304316 69028
rect 304816 69080 304868 69086
rect 304816 69022 304868 69028
rect 303540 6798 303568 69022
rect 304356 9512 304408 9518
rect 304356 9454 304408 9460
rect 303528 6792 303580 6798
rect 303528 6734 303580 6740
rect 303436 6724 303488 6730
rect 303436 6666 303488 6672
rect 304368 480 304396 9454
rect 304828 6662 304856 69022
rect 304816 6656 304868 6662
rect 304816 6598 304868 6604
rect 304920 6594 304948 71726
rect 305656 69086 305684 71726
rect 306300 71726 306337 71754
rect 307007 71754 307035 72012
rect 307705 71754 307733 72012
rect 307007 71726 307064 71754
rect 305644 69080 305696 69086
rect 305644 69022 305696 69028
rect 306196 69080 306248 69086
rect 306196 69022 306248 69028
rect 304908 6588 304960 6594
rect 304908 6530 304960 6536
rect 306208 6526 306236 69022
rect 306196 6520 306248 6526
rect 306196 6462 306248 6468
rect 306300 6458 306328 71726
rect 307036 69086 307064 71726
rect 307588 71726 307733 71754
rect 308403 71754 308431 72012
rect 309101 71754 309129 72012
rect 309798 71754 309826 72012
rect 308403 71726 308444 71754
rect 307024 69080 307076 69086
rect 307024 69022 307076 69028
rect 306380 13524 306432 13530
rect 306380 13466 306432 13472
rect 306288 6452 306340 6458
rect 306288 6394 306340 6400
rect 305552 2916 305604 2922
rect 305552 2858 305604 2864
rect 305564 480 305592 2858
rect 306392 490 306420 13466
rect 307588 6322 307616 71726
rect 308416 69086 308444 71726
rect 308968 71726 309129 71754
rect 309796 71726 309826 71754
rect 310496 71754 310524 72012
rect 311194 71754 311222 72012
rect 310496 71726 310560 71754
rect 307668 69080 307720 69086
rect 307668 69022 307720 69028
rect 308404 69080 308456 69086
rect 308404 69022 308456 69028
rect 307680 6390 307708 69022
rect 308968 9654 308996 71726
rect 309796 69086 309824 71726
rect 310152 69624 310204 69630
rect 310152 69566 310204 69572
rect 309876 69284 309928 69290
rect 309876 69226 309928 69232
rect 309048 69080 309100 69086
rect 309048 69022 309100 69028
rect 309784 69080 309836 69086
rect 309784 69022 309836 69028
rect 308956 9648 309008 9654
rect 308956 9590 309008 9596
rect 307944 9308 307996 9314
rect 307944 9250 307996 9256
rect 307668 6384 307720 6390
rect 307668 6326 307720 6332
rect 307576 6316 307628 6322
rect 307576 6258 307628 6264
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 9250
rect 309060 6254 309088 69022
rect 309888 64874 309916 69226
rect 310164 67182 310192 69566
rect 310336 69420 310388 69426
rect 310336 69362 310388 69368
rect 310348 68678 310376 69362
rect 310532 69154 310560 71726
rect 311176 71726 311222 71754
rect 311892 71754 311920 72012
rect 312590 71754 312618 72012
rect 311892 71726 311940 71754
rect 310520 69148 310572 69154
rect 310520 69090 310572 69096
rect 311176 69086 311204 71726
rect 311808 69148 311860 69154
rect 311808 69090 311860 69096
rect 310428 69080 310480 69086
rect 310428 69022 310480 69028
rect 311164 69080 311216 69086
rect 311164 69022 311216 69028
rect 311716 69080 311768 69086
rect 311716 69022 311768 69028
rect 310336 68672 310388 68678
rect 310336 68614 310388 68620
rect 310152 67176 310204 67182
rect 310152 67118 310204 67124
rect 309796 64846 309916 64874
rect 309796 15978 309824 64846
rect 309784 15972 309836 15978
rect 309784 15914 309836 15920
rect 309784 14748 309836 14754
rect 309784 14690 309836 14696
rect 309048 6248 309100 6254
rect 309048 6190 309100 6196
rect 309048 2848 309100 2854
rect 309048 2790 309100 2796
rect 309060 480 309088 2790
rect 309796 490 309824 14690
rect 310440 6186 310468 69022
rect 311728 9314 311756 69022
rect 311820 9518 311848 69090
rect 311912 69086 311940 71726
rect 312556 71726 312618 71754
rect 313287 71754 313315 72012
rect 313985 71754 314013 72012
rect 313287 71726 313320 71754
rect 311900 69080 311952 69086
rect 311900 69022 311952 69028
rect 312556 68610 312584 71726
rect 313188 69624 313240 69630
rect 313188 69566 313240 69572
rect 313096 69080 313148 69086
rect 313096 69022 313148 69028
rect 312544 68604 312596 68610
rect 312544 68546 312596 68552
rect 311808 9512 311860 9518
rect 311808 9454 311860 9460
rect 311716 9308 311768 9314
rect 311716 9250 311768 9256
rect 313108 9246 313136 69022
rect 311440 9240 311492 9246
rect 311440 9182 311492 9188
rect 313096 9240 313148 9246
rect 313096 9182 313148 9188
rect 310428 6180 310480 6186
rect 310428 6122 310480 6128
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 9182
rect 313200 3602 313228 69566
rect 313292 18630 313320 71726
rect 313476 71726 314013 71754
rect 314683 71754 314711 72012
rect 315381 71754 315409 72012
rect 316079 71754 316107 72012
rect 316776 71754 316804 72012
rect 314683 71726 314884 71754
rect 313280 18624 313332 18630
rect 313280 18566 313332 18572
rect 313476 16114 313504 71726
rect 314752 68604 314804 68610
rect 314752 68546 314804 68552
rect 313464 16108 313516 16114
rect 313464 16050 313516 16056
rect 313832 12232 313884 12238
rect 313832 12174 313884 12180
rect 312636 3596 312688 3602
rect 312636 3538 312688 3544
rect 313188 3596 313240 3602
rect 313188 3538 313240 3544
rect 312648 480 312676 3538
rect 313844 480 313872 12174
rect 314764 3505 314792 68546
rect 314750 3496 314806 3505
rect 314750 3431 314806 3440
rect 314856 3369 314884 71726
rect 315316 71726 315409 71754
rect 316052 71726 316107 71754
rect 316420 71726 316804 71754
rect 317474 71754 317502 72012
rect 318172 71754 318200 72012
rect 317474 71726 317552 71754
rect 315316 68610 315344 71726
rect 315304 68604 315356 68610
rect 315304 68546 315356 68552
rect 315028 8424 315080 8430
rect 315028 8366 315080 8372
rect 314842 3360 314898 3369
rect 314842 3295 314898 3304
rect 315040 480 315068 8366
rect 316052 3466 316080 71726
rect 316316 16040 316368 16046
rect 316316 15982 316368 15988
rect 316224 3596 316276 3602
rect 316224 3538 316276 3544
rect 316040 3460 316092 3466
rect 316040 3402 316092 3408
rect 316236 480 316264 3538
rect 316328 3346 316356 15982
rect 316420 3534 316448 71726
rect 317524 3670 317552 71726
rect 317616 71726 318200 71754
rect 318870 71754 318898 72012
rect 319568 71754 319596 72012
rect 318870 71726 318932 71754
rect 317512 3664 317564 3670
rect 317512 3606 317564 3612
rect 316408 3528 316460 3534
rect 316408 3470 316460 3476
rect 317616 3466 317644 71726
rect 318524 8492 318576 8498
rect 318524 8434 318576 8440
rect 317604 3460 317656 3466
rect 317604 3402 317656 3408
rect 316328 3318 317368 3346
rect 317340 480 317368 3318
rect 318536 480 318564 8434
rect 318904 3738 318932 71726
rect 319548 71726 319596 71754
rect 320265 71754 320293 72012
rect 320963 71754 320991 72012
rect 320265 71726 320312 71754
rect 319548 69290 319576 71726
rect 320284 69494 320312 71726
rect 320376 71726 320991 71754
rect 321560 71800 321612 71806
rect 321560 71742 321612 71748
rect 321661 71754 321689 72012
rect 322359 71806 322387 72012
rect 322347 71800 322399 71806
rect 320272 69488 320324 69494
rect 320272 69430 320324 69436
rect 319536 69284 319588 69290
rect 319536 69226 319588 69232
rect 320180 68808 320232 68814
rect 320180 68750 320232 68756
rect 320192 16574 320220 68750
rect 320376 17338 320404 71726
rect 320364 17332 320416 17338
rect 320364 17274 320416 17280
rect 320192 16546 320496 16574
rect 318892 3732 318944 3738
rect 318892 3674 318944 3680
rect 319720 3664 319772 3670
rect 319720 3606 319772 3612
rect 319732 480 319760 3606
rect 320468 490 320496 16546
rect 321572 14822 321600 71742
rect 321661 71726 321692 71754
rect 323057 71754 323085 72012
rect 323754 71754 323782 72012
rect 322347 71742 322399 71748
rect 321664 17270 321692 71726
rect 323044 71726 323085 71754
rect 323136 71726 323782 71754
rect 324320 71800 324372 71806
rect 324452 71754 324480 72012
rect 325150 71806 325178 72012
rect 324320 71742 324372 71748
rect 323044 69562 323072 71726
rect 323032 69556 323084 69562
rect 323032 69498 323084 69504
rect 321652 17264 321704 17270
rect 321652 17206 321704 17212
rect 323136 16182 323164 71726
rect 324228 69556 324280 69562
rect 324228 69498 324280 69504
rect 323124 16176 323176 16182
rect 323124 16118 323176 16124
rect 321560 14816 321612 14822
rect 321560 14758 321612 14764
rect 322112 8560 322164 8566
rect 322112 8502 322164 8508
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 8502
rect 324240 3534 324268 69498
rect 324332 14890 324360 71742
rect 324424 71726 324480 71754
rect 325138 71800 325190 71806
rect 325848 71754 325876 72012
rect 326546 71754 326574 72012
rect 325138 71742 325190 71748
rect 325804 71726 325876 71754
rect 326540 71726 326574 71754
rect 327080 71800 327132 71806
rect 327243 71754 327271 72012
rect 327941 71806 327969 72012
rect 327080 71742 327132 71748
rect 324424 17406 324452 71726
rect 325804 70310 325832 71726
rect 325792 70304 325844 70310
rect 325792 70246 325844 70252
rect 326540 67250 326568 71726
rect 326528 67244 326580 67250
rect 326528 67186 326580 67192
rect 324412 17400 324464 17406
rect 324412 17342 324464 17348
rect 327092 16250 327120 71742
rect 327184 71726 327271 71754
rect 327929 71800 327981 71806
rect 327929 71742 327981 71748
rect 328460 71800 328512 71806
rect 328639 71754 328667 72012
rect 329337 71806 329365 72012
rect 328460 71742 328512 71748
rect 327184 18698 327212 71726
rect 327724 69148 327776 69154
rect 327724 69090 327776 69096
rect 327172 18692 327224 18698
rect 327172 18634 327224 18640
rect 327080 16244 327132 16250
rect 327080 16186 327132 16192
rect 324320 14884 324372 14890
rect 324320 14826 324372 14832
rect 327736 13598 327764 69090
rect 328472 17474 328500 71742
rect 328564 71726 328667 71754
rect 329325 71800 329377 71806
rect 329325 71742 329377 71748
rect 329840 71800 329892 71806
rect 330035 71754 330063 72012
rect 330732 71806 330760 72012
rect 329840 71742 329892 71748
rect 328564 44878 328592 71726
rect 328552 44872 328604 44878
rect 328552 44814 328604 44820
rect 329852 18766 329880 71742
rect 329944 71726 330063 71754
rect 330720 71800 330772 71806
rect 330720 71742 330772 71748
rect 331220 71800 331272 71806
rect 331430 71754 331458 72012
rect 332128 71806 332156 72012
rect 331220 71742 331272 71748
rect 329944 22778 329972 71726
rect 329932 22772 329984 22778
rect 329932 22714 329984 22720
rect 329840 18760 329892 18766
rect 329840 18702 329892 18708
rect 328460 17468 328512 17474
rect 328460 17410 328512 17416
rect 331232 14958 331260 71742
rect 331416 71726 331458 71754
rect 332116 71800 332168 71806
rect 332826 71754 332854 72012
rect 332116 71742 332168 71748
rect 332796 71726 332854 71754
rect 333524 71754 333552 72012
rect 333980 71800 334032 71806
rect 333524 71726 333560 71754
rect 334221 71754 334249 72012
rect 334919 71806 334947 72012
rect 333980 71742 334032 71748
rect 331312 47592 331364 47598
rect 331312 47534 331364 47540
rect 331324 16574 331352 47534
rect 331416 25566 331444 71726
rect 332796 69154 332824 71726
rect 332784 69148 332836 69154
rect 332784 69090 332836 69096
rect 333532 69086 333560 71726
rect 331864 69080 331916 69086
rect 331864 69022 331916 69028
rect 333520 69080 333572 69086
rect 333520 69022 333572 69028
rect 331876 50386 331904 69022
rect 331864 50380 331916 50386
rect 331864 50322 331916 50328
rect 331404 25560 331456 25566
rect 331404 25502 331456 25508
rect 331324 16546 331628 16574
rect 331220 14952 331272 14958
rect 331220 14894 331272 14900
rect 327724 13592 327776 13598
rect 327724 13534 327776 13540
rect 324412 13456 324464 13462
rect 324412 13398 324464 13404
rect 323308 3528 323360 3534
rect 323308 3470 323360 3476
rect 324228 3528 324280 3534
rect 324228 3470 324280 3476
rect 323320 480 323348 3470
rect 324424 480 324452 13398
rect 328000 13388 328052 13394
rect 328000 13330 328052 13336
rect 325608 8628 325660 8634
rect 325608 8570 325660 8576
rect 325620 480 325648 8570
rect 326804 3596 326856 3602
rect 326804 3538 326856 3544
rect 326816 480 326844 3538
rect 328012 480 328040 13330
rect 329196 8696 329248 8702
rect 329196 8638 329248 8644
rect 329208 480 329236 8638
rect 330392 3664 330444 3670
rect 330392 3606 330444 3612
rect 330404 480 330432 3606
rect 331600 480 331628 16546
rect 332692 8764 332744 8770
rect 332692 8706 332744 8712
rect 332704 480 332732 8706
rect 333888 3732 333940 3738
rect 333888 3674 333940 3680
rect 333900 480 333928 3674
rect 333992 3641 334020 71742
rect 334084 71726 334249 71754
rect 334907 71800 334959 71806
rect 334907 71742 334959 71748
rect 335452 71800 335504 71806
rect 335617 71754 335645 72012
rect 336315 71806 336343 72012
rect 335452 71742 335504 71748
rect 334084 17610 334112 71726
rect 334072 17604 334124 17610
rect 334072 17546 334124 17552
rect 334624 14680 334676 14686
rect 334624 14622 334676 14628
rect 333978 3632 334034 3641
rect 333978 3567 334034 3576
rect 334636 490 334664 14622
rect 335464 3806 335492 71742
rect 335556 71726 335645 71754
rect 336303 71800 336355 71806
rect 337013 71754 337041 72012
rect 337710 71754 337738 72012
rect 336303 71742 336355 71748
rect 336752 71726 337041 71754
rect 337120 71726 337738 71754
rect 338120 71800 338172 71806
rect 338120 71742 338172 71748
rect 335452 3800 335504 3806
rect 335556 3777 335584 71726
rect 336280 8832 336332 8838
rect 336280 8774 336332 8780
rect 335452 3742 335504 3748
rect 335542 3768 335598 3777
rect 335542 3703 335598 3712
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 8774
rect 336752 3874 336780 71726
rect 337120 64874 337148 71726
rect 338028 70304 338080 70310
rect 338028 70246 338080 70252
rect 336844 64846 337148 64874
rect 336844 3942 336872 64846
rect 336832 3936 336884 3942
rect 336832 3878 336884 3884
rect 336740 3868 336792 3874
rect 336740 3810 336792 3816
rect 338040 3330 338068 70246
rect 338132 4078 338160 71742
rect 338304 49020 338356 49026
rect 338304 48962 338356 48968
rect 338120 4072 338172 4078
rect 338120 4014 338172 4020
rect 338316 3482 338344 48962
rect 338408 4010 338436 72012
rect 339106 71806 339134 72012
rect 339094 71800 339146 71806
rect 339804 71754 339832 72012
rect 340502 71754 340530 72012
rect 339094 71742 339146 71748
rect 339604 71726 339832 71754
rect 339880 71726 340530 71754
rect 340972 71800 341024 71806
rect 341199 71754 341227 72012
rect 341897 71806 341925 72012
rect 342595 71890 342623 72012
rect 342364 71862 342623 71890
rect 340972 71742 341024 71748
rect 339604 4146 339632 71726
rect 339880 64874 339908 71726
rect 339696 64846 339908 64874
rect 339592 4140 339644 4146
rect 339592 4082 339644 4088
rect 338396 4004 338448 4010
rect 338396 3946 338448 3952
rect 338316 3454 338712 3482
rect 337476 3324 337528 3330
rect 337476 3266 337528 3272
rect 338028 3324 338080 3330
rect 338028 3266 338080 3272
rect 337488 480 337516 3266
rect 338684 480 338712 3454
rect 339696 3398 339724 64846
rect 339868 8900 339920 8906
rect 339868 8842 339920 8848
rect 339684 3392 339736 3398
rect 339684 3334 339736 3340
rect 339880 480 339908 8842
rect 340984 3874 341012 71742
rect 341168 71726 341227 71754
rect 341885 71800 341937 71806
rect 341885 71742 341937 71748
rect 341064 11960 341116 11966
rect 341064 11902 341116 11908
rect 340972 3868 341024 3874
rect 340972 3810 341024 3816
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 340984 480 341012 3334
rect 341076 3074 341104 11902
rect 341168 3194 341196 71726
rect 342364 70174 342392 71862
rect 343293 71754 343321 72012
rect 343991 71754 344019 72012
rect 344688 71754 344716 72012
rect 342456 71726 343321 71754
rect 343652 71726 344019 71754
rect 344204 71726 344716 71754
rect 345386 71754 345414 72012
rect 346084 71754 346112 72012
rect 346782 71754 346810 72012
rect 347480 71754 347508 72012
rect 348177 71754 348205 72012
rect 345386 71726 345428 71754
rect 342352 70168 342404 70174
rect 342352 70110 342404 70116
rect 342168 69488 342220 69494
rect 342168 69430 342220 69436
rect 342180 3398 342208 69430
rect 342352 19984 342404 19990
rect 342352 19926 342404 19932
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 341156 3188 341208 3194
rect 341156 3130 341208 3136
rect 341076 3046 342208 3074
rect 342180 480 342208 3046
rect 342364 626 342392 19926
rect 342456 3126 342484 71726
rect 342444 3120 342496 3126
rect 342444 3062 342496 3068
rect 343652 3058 343680 71726
rect 344204 64874 344232 71726
rect 345400 70242 345428 71726
rect 346044 71726 346112 71754
rect 346412 71726 346810 71754
rect 347424 71726 347508 71754
rect 347976 71726 348205 71754
rect 348875 71754 348903 72012
rect 349252 71800 349304 71806
rect 348875 71726 348924 71754
rect 349573 71754 349601 72012
rect 350271 71806 350299 72012
rect 350969 71890 350997 72012
rect 350644 71862 350997 71890
rect 349252 71742 349304 71748
rect 346044 70378 346072 71726
rect 346032 70372 346084 70378
rect 346032 70314 346084 70320
rect 345388 70236 345440 70242
rect 345388 70178 345440 70184
rect 345020 68740 345072 68746
rect 345020 68682 345072 68688
rect 343744 64846 344232 64874
rect 343744 3806 343772 64846
rect 345032 16574 345060 68682
rect 345032 16546 345336 16574
rect 344560 4004 344612 4010
rect 344560 3946 344612 3952
rect 343732 3800 343784 3806
rect 343732 3742 343784 3748
rect 343640 3052 343692 3058
rect 343640 2994 343692 3000
rect 342364 598 342944 626
rect 342916 490 342944 598
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
<<<<<<< HEAD
rect 343334 -960 343446 480
rect 344530 -960 344642 480
=======
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3946
rect 345308 490 345336 16546
rect 346412 2922 346440 71726
rect 347424 64874 347452 71726
rect 346504 64846 347452 64874
rect 346504 3398 346532 64846
rect 346952 12436 347004 12442
rect 346952 12378 347004 12384
rect 346492 3392 346544 3398
rect 346492 3334 346544 3340
rect 346400 2916 346452 2922
rect 346400 2858 346452 2864
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 12378
rect 347976 2854 348004 71726
rect 348896 69630 348924 71726
rect 348884 69624 348936 69630
rect 348884 69566 348936 69572
rect 349264 16574 349292 71742
rect 349172 16546 349292 16574
rect 349448 71726 349601 71754
rect 350259 71800 350311 71806
rect 350259 71742 350311 71748
rect 348056 3596 348108 3602
rect 348056 3538 348108 3544
rect 347964 2848 348016 2854
rect 347964 2790 348016 2796
rect 348068 480 348096 3538
rect 349172 3534 349200 16546
rect 349344 15020 349396 15026
rect 349344 14962 349396 14968
rect 349252 13320 349304 13326
rect 349252 13262 349304 13268
rect 349160 3528 349212 3534
rect 349160 3470 349212 3476
rect 349264 480 349292 13262
rect 349356 3346 349384 14962
rect 349448 3466 349476 71726
rect 350644 69562 350672 71862
rect 351666 71754 351694 72012
rect 352364 71754 352392 72012
rect 353062 71754 353090 72012
rect 350736 71726 351694 71754
rect 351932 71726 352392 71754
rect 352484 71726 353090 71754
rect 353760 71754 353788 72012
rect 354458 71754 354486 72012
rect 355155 71754 355183 72012
rect 355853 71754 355881 72012
rect 356551 71754 356579 72012
rect 357249 71754 357277 72012
rect 357947 71754 357975 72012
rect 353760 71726 353800 71754
rect 350632 69556 350684 69562
rect 350632 69498 350684 69504
rect 350736 3670 350764 71726
rect 351932 3806 351960 71726
rect 352484 64874 352512 71726
rect 353772 70310 353800 71726
rect 354416 71726 354486 71754
rect 354692 71726 355183 71754
rect 355244 71726 355881 71754
rect 356164 71726 356579 71754
rect 356992 71726 357277 71754
rect 357452 71726 357975 71754
rect 358644 71754 358672 72012
rect 359342 71754 359370 72012
rect 360040 71754 360068 72012
rect 358644 71726 358768 71754
rect 359342 71726 359412 71754
rect 353760 70304 353812 70310
rect 353760 70246 353812 70252
rect 353944 69964 353996 69970
rect 353944 69906 353996 69912
rect 352024 64846 352512 64874
rect 352024 3942 352052 64846
rect 352840 14612 352892 14618
rect 352840 14554 352892 14560
rect 352012 3936 352064 3942
rect 352012 3878 352064 3884
rect 351920 3800 351972 3806
rect 351920 3742 351972 3748
rect 350724 3664 350776 3670
rect 350724 3606 350776 3612
rect 349436 3460 349488 3466
rect 349436 3402 349488 3408
rect 349356 3318 350488 3346
rect 350460 480 350488 3318
rect 351644 2984 351696 2990
rect 351644 2926 351696 2932
rect 351656 480 351684 2926
rect 352852 480 352880 14554
rect 353956 11966 353984 69906
rect 354416 69494 354444 71726
rect 354404 69488 354456 69494
rect 354404 69430 354456 69436
rect 354036 21412 354088 21418
rect 354036 21354 354088 21360
rect 353944 11960 353996 11966
rect 353944 11902 353996 11908
rect 354048 6914 354076 21354
rect 354128 16380 354180 16386
rect 354128 16322 354180 16328
rect 353956 6886 354076 6914
rect 353956 3670 353984 6886
rect 354036 4276 354088 4282
rect 354036 4218 354088 4224
rect 353944 3664 353996 3670
rect 353944 3606 353996 3612
rect 354048 480 354076 4218
rect 354140 3466 354168 16322
rect 354692 4010 354720 71726
rect 355244 64874 355272 71726
rect 354784 64846 355272 64874
rect 354680 4004 354732 4010
rect 354680 3946 354732 3952
rect 354784 3602 354812 64846
rect 354772 3596 354824 3602
rect 354772 3538 354824 3544
rect 355232 3528 355284 3534
rect 355232 3470 355284 3476
rect 354128 3460 354180 3466
rect 354128 3402 354180 3408
rect 355244 480 355272 3470
rect 356164 2990 356192 71726
rect 356992 64874 357020 71726
rect 356256 64846 357020 64874
rect 356256 3534 356284 64846
rect 356336 7064 356388 7070
rect 356336 7006 356388 7012
rect 356244 3528 356296 3534
rect 356244 3470 356296 3476
rect 356152 2984 356204 2990
rect 356152 2926 356204 2932
rect 356348 480 356376 7006
rect 357452 3534 357480 71726
rect 358740 6914 358768 71726
rect 359384 69086 359412 71726
rect 360028 71726 360068 71754
rect 360738 71754 360766 72012
rect 361436 71754 361464 72012
rect 362133 71754 362161 72012
rect 362831 71754 362859 72012
rect 363529 71754 363557 72012
rect 364227 71754 364255 72012
rect 364925 71754 364953 72012
rect 365622 71754 365650 72012
rect 360738 71726 360792 71754
rect 361436 71726 361528 71754
rect 362133 71726 362172 71754
rect 359372 69080 359424 69086
rect 359372 69022 359424 69028
rect 359924 7132 359976 7138
rect 359924 7074 359976 7080
rect 358648 6886 358768 6914
rect 357532 3664 357584 3670
rect 357532 3606 357584 3612
rect 357440 3528 357492 3534
rect 357440 3470 357492 3476
rect 357544 480 357572 3606
rect 358648 3602 358676 6886
rect 358636 3596 358688 3602
rect 358636 3538 358688 3544
rect 358728 3528 358780 3534
rect 358728 3470 358780 3476
rect 358740 480 358768 3470
rect 359936 480 359964 7074
rect 360028 3670 360056 71726
rect 360764 69086 360792 71726
rect 360108 69080 360160 69086
rect 360108 69022 360160 69028
rect 360752 69080 360804 69086
rect 360752 69022 360804 69028
rect 361396 69080 361448 69086
rect 361396 69022 361448 69028
rect 360016 3664 360068 3670
rect 360016 3606 360068 3612
rect 360120 3194 360148 69022
rect 360844 13728 360896 13734
rect 360844 13670 360896 13676
rect 360856 3942 360884 13670
rect 361408 4146 361436 69022
rect 361396 4140 361448 4146
rect 361396 4082 361448 4088
rect 361500 4010 361528 71726
rect 362144 69086 362172 71726
rect 362788 71726 362859 71754
rect 363524 71726 363557 71754
rect 364168 71726 364255 71754
rect 364904 71726 364953 71754
rect 365548 71726 365650 71754
rect 366320 71754 366348 72012
rect 367018 71754 367046 72012
rect 367716 71754 367744 72012
rect 368414 71754 368442 72012
rect 366320 71726 366404 71754
rect 367018 71726 367048 71754
rect 367716 71726 367784 71754
rect 362132 69080 362184 69086
rect 362132 69022 362184 69028
rect 361488 4004 361540 4010
rect 361488 3946 361540 3952
rect 360844 3936 360896 3942
rect 360844 3878 360896 3884
rect 362788 3806 362816 71726
rect 363524 69086 363552 71726
rect 362868 69080 362920 69086
rect 362868 69022 362920 69028
rect 363512 69080 363564 69086
rect 363512 69022 363564 69028
rect 362880 3874 362908 69022
rect 363512 7200 363564 7206
rect 363512 7142 363564 7148
rect 362868 3868 362920 3874
rect 362868 3810 362920 3816
rect 362776 3800 362828 3806
rect 362776 3742 362828 3748
rect 362316 3596 362368 3602
rect 362316 3538 362368 3544
rect 361120 3460 361172 3466
rect 361120 3402 361172 3408
rect 360108 3188 360160 3194
rect 360108 3130 360160 3136
rect 361132 480 361160 3402
rect 362328 480 362356 3538
rect 363524 480 363552 7142
rect 364168 3670 364196 71726
rect 364904 69086 364932 71726
rect 364248 69080 364300 69086
rect 364248 69022 364300 69028
rect 364892 69080 364944 69086
rect 364892 69022 364944 69028
rect 364260 3738 364288 69022
rect 364616 3936 364668 3942
rect 364616 3878 364668 3884
rect 364248 3732 364300 3738
rect 364248 3674 364300 3680
rect 364156 3664 364208 3670
rect 364156 3606 364208 3612
rect 364628 480 364656 3878
rect 365548 3466 365576 71726
rect 366376 69086 366404 71726
rect 365628 69080 365680 69086
rect 365628 69022 365680 69028
rect 366364 69080 366416 69086
rect 366364 69022 366416 69028
rect 366916 69080 366968 69086
rect 366916 69022 366968 69028
rect 365640 3534 365668 69022
rect 366928 16574 366956 69022
rect 366836 16546 366956 16574
rect 365628 3528 365680 3534
rect 365628 3470 365680 3476
rect 365536 3460 365588 3466
rect 365536 3402 365588 3408
rect 366836 3330 366864 16546
rect 367020 11778 367048 71726
rect 367756 69426 367784 71726
rect 368400 71726 368442 71754
rect 369111 71754 369139 72012
rect 369809 71754 369837 72012
rect 369111 71726 369164 71754
rect 367744 69420 367796 69426
rect 367744 69362 367796 69368
rect 367100 17536 367152 17542
rect 367100 17478 367152 17484
rect 367112 16574 367140 17478
rect 367112 16546 367784 16574
rect 366928 11750 367048 11778
rect 366824 3324 366876 3330
rect 366824 3266 366876 3272
rect 365812 3188 365864 3194
rect 365812 3130 365864 3136
rect 365824 480 365852 3130
rect 366928 2854 366956 11750
rect 367008 7268 367060 7274
rect 367008 7210 367060 7216
rect 366916 2848 366968 2854
rect 366916 2790 366968 2796
rect 367020 480 367048 7210
rect 367756 490 367784 16546
rect 368400 2922 368428 71726
rect 369136 69086 369164 71726
rect 369780 71726 369837 71754
rect 370507 71754 370535 72012
rect 371205 71754 371233 72012
rect 371903 71754 371931 72012
rect 370507 71726 370544 71754
rect 369124 69080 369176 69086
rect 369124 69022 369176 69028
rect 369676 69080 369728 69086
rect 369676 69022 369728 69028
rect 369400 3596 369452 3602
rect 369400 3538 369452 3544
rect 368388 2916 368440 2922
rect 368388 2858 368440 2864
rect 368032 598 368244 626
rect 368032 490 368060 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
<<<<<<< HEAD
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
=======
rect 367756 462 368060 490
rect 368216 480 368244 598
rect 369412 480 369440 3538
rect 369688 2990 369716 69022
rect 369780 3058 369808 71726
rect 370516 69494 370544 71726
rect 371160 71726 371233 71754
rect 371896 71726 371931 71754
rect 372600 71754 372628 72012
rect 373298 71754 373326 72012
rect 372600 71726 372660 71754
rect 370504 69488 370556 69494
rect 370504 69430 370556 69436
rect 370596 7336 370648 7342
rect 370596 7278 370648 7284
rect 369768 3052 369820 3058
rect 369768 2994 369820 3000
rect 369676 2984 369728 2990
rect 369676 2926 369728 2932
rect 370608 480 370636 7278
rect 371160 3126 371188 71726
rect 371792 69896 371844 69902
rect 371792 69838 371844 69844
rect 371804 64874 371832 69838
rect 371896 69562 371924 71726
rect 372632 69630 372660 71726
rect 373276 71726 373326 71754
rect 373996 71754 374024 72012
rect 374694 71754 374722 72012
rect 373996 71726 374040 71754
rect 374694 71726 374776 71754
rect 372620 69624 372672 69630
rect 372620 69566 372672 69572
rect 371884 69556 371936 69562
rect 371884 69498 371936 69504
rect 373276 69086 373304 71726
rect 374012 70378 374040 71726
rect 374000 70372 374052 70378
rect 374000 70314 374052 70320
rect 374748 69086 374776 71726
rect 375392 70310 375420 72012
rect 376089 71754 376117 72012
rect 376787 71754 376815 72012
rect 376089 71726 376156 71754
rect 375380 70304 375432 70310
rect 375380 70246 375432 70252
rect 376128 69086 376156 71726
rect 376772 71726 376815 71754
rect 377485 71754 377513 72012
rect 378183 71754 378211 72012
rect 378881 71754 378909 72012
rect 379578 71754 379606 72012
rect 380276 71754 380304 72012
rect 377485 71726 377536 71754
rect 378183 71726 378272 71754
rect 378881 71726 378916 71754
rect 379578 71726 379652 71754
rect 376772 69358 376800 71726
rect 376760 69352 376812 69358
rect 376760 69294 376812 69300
rect 377508 69086 377536 71726
rect 378244 70174 378272 71726
rect 378232 70168 378284 70174
rect 378232 70110 378284 70116
rect 378888 69086 378916 71726
rect 379624 70242 379652 71726
rect 380268 71726 380304 71754
rect 380974 71754 381002 72012
rect 381672 71754 381700 72012
rect 380974 71726 381032 71754
rect 379612 70236 379664 70242
rect 379612 70178 379664 70184
rect 380268 69086 380296 71726
rect 381004 69970 381032 71726
rect 381648 71726 381700 71754
rect 382370 71754 382398 72012
rect 383067 71754 383095 72012
rect 383765 71754 383793 72012
rect 382370 71726 382412 71754
rect 383067 71726 383516 71754
rect 380992 69964 381044 69970
rect 380992 69906 381044 69912
rect 381648 69086 381676 71726
rect 382384 69086 382412 71726
rect 373264 69080 373316 69086
rect 373264 69022 373316 69028
rect 373908 69080 373960 69086
rect 373908 69022 373960 69028
rect 374736 69080 374788 69086
rect 374736 69022 374788 69028
rect 375288 69080 375340 69086
rect 375288 69022 375340 69028
rect 376116 69080 376168 69086
rect 376116 69022 376168 69028
rect 376668 69080 376720 69086
rect 376668 69022 376720 69028
rect 377496 69080 377548 69086
rect 377496 69022 377548 69028
rect 378048 69080 378100 69086
rect 378048 69022 378100 69028
rect 378876 69080 378928 69086
rect 378876 69022 378928 69028
rect 379428 69080 379480 69086
rect 379428 69022 379480 69028
rect 380256 69080 380308 69086
rect 380256 69022 380308 69028
rect 380808 69080 380860 69086
rect 380808 69022 380860 69028
rect 381636 69080 381688 69086
rect 381636 69022 381688 69028
rect 382188 69080 382240 69086
rect 382188 69022 382240 69028
rect 382372 69080 382424 69086
rect 382372 69022 382424 69028
rect 371804 64846 371924 64874
rect 371240 16312 371292 16318
rect 371240 16254 371292 16260
rect 371148 3120 371200 3126
rect 371148 3062 371200 3068
rect 371252 490 371280 16254
rect 371896 7342 371924 64846
rect 371884 7336 371936 7342
rect 371884 7278 371936 7284
rect 372896 4140 372948 4146
rect 372896 4082 372948 4088
rect 371528 598 371740 626
rect 371528 490 371556 598
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 462 371556 490
rect 371712 480 371740 598
rect 372908 480 372936 4082
rect 373920 3194 373948 69022
rect 374000 67312 374052 67318
rect 374000 67254 374052 67260
rect 374012 3262 374040 67254
rect 374092 7404 374144 7410
rect 374092 7346 374144 7352
rect 374000 3256 374052 3262
rect 374000 3198 374052 3204
rect 373908 3188 373960 3194
rect 373908 3130 373960 3136
rect 374104 480 374132 7346
rect 375300 6914 375328 69022
rect 375208 6886 375328 6914
rect 375208 3330 375236 6886
rect 376484 4004 376536 4010
rect 376484 3946 376536 3952
rect 375196 3324 375248 3330
rect 375196 3266 375248 3272
rect 375288 3256 375340 3262
rect 375288 3198 375340 3204
rect 375300 480 375328 3198
rect 376496 480 376524 3946
rect 376680 3330 376708 69022
rect 377680 7472 377732 7478
rect 377680 7414 377732 7420
rect 376668 3324 376720 3330
rect 376668 3266 376720 3272
rect 377692 480 377720 7414
rect 378060 3398 378088 69022
rect 378416 9784 378468 9790
rect 378416 9726 378468 9732
rect 378048 3392 378100 3398
rect 378048 3334 378100 3340
rect 378428 490 378456 9726
rect 379440 4146 379468 69022
rect 379428 4140 379480 4146
rect 379428 4082 379480 4088
rect 380820 4078 380848 69022
rect 381176 7540 381228 7546
rect 381176 7482 381228 7488
rect 380808 4072 380860 4078
rect 380808 4014 380860 4020
rect 379980 3868 380032 3874
rect 379980 3810 380032 3816
rect 378704 598 378916 626
rect 378704 490 378732 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 3810
rect 381188 480 381216 7482
rect 382200 4010 382228 69022
rect 383488 64394 383516 71726
rect 383764 71726 383793 71754
rect 384463 71754 384491 72012
rect 385161 71754 385189 72012
rect 384463 71726 384528 71754
rect 383764 69290 383792 71726
rect 383752 69284 383804 69290
rect 383752 69226 383804 69232
rect 383568 69080 383620 69086
rect 383568 69022 383620 69028
rect 383476 64388 383528 64394
rect 383476 64330 383528 64336
rect 383580 17270 383608 69022
rect 384500 68882 384528 71726
rect 385144 71726 385189 71754
rect 385859 71754 385887 72012
rect 386556 71754 386584 72012
rect 387254 71754 387282 72012
rect 387952 71754 387980 72012
rect 388650 71754 388678 72012
rect 385859 71726 385908 71754
rect 386556 71726 386644 71754
rect 387254 71726 387288 71754
rect 387952 71726 388024 71754
rect 384488 68876 384540 68882
rect 384488 68818 384540 68824
rect 385144 67318 385172 71726
rect 385880 69086 385908 71726
rect 385868 69080 385920 69086
rect 385868 69022 385920 69028
rect 386328 69080 386380 69086
rect 386328 69022 386380 69028
rect 385132 67312 385184 67318
rect 385132 67254 385184 67260
rect 386340 18630 386368 69022
rect 386616 68814 386644 71726
rect 386604 68808 386656 68814
rect 386604 68750 386656 68756
rect 387260 67250 387288 71726
rect 387248 67244 387300 67250
rect 387248 67186 387300 67192
rect 387996 65890 388024 71726
rect 388640 71726 388678 71754
rect 389348 71754 389376 72012
rect 390045 71754 390073 72012
rect 389348 71726 389404 71754
rect 388640 69086 388668 71726
rect 389376 69154 389404 71726
rect 390020 71726 390073 71754
rect 390743 71754 390771 72012
rect 391441 71754 391469 72012
rect 392139 71754 392167 72012
rect 390743 71726 390784 71754
rect 391441 71726 391520 71754
rect 389364 69148 389416 69154
rect 389364 69090 389416 69096
rect 390020 69086 390048 71726
rect 390376 69148 390428 69154
rect 390376 69090 390428 69096
rect 388628 69080 388680 69086
rect 388628 69022 388680 69028
rect 389088 69080 389140 69086
rect 389088 69022 389140 69028
rect 390008 69080 390060 69086
rect 390008 69022 390060 69028
rect 387984 65884 388036 65890
rect 387984 65826 388036 65832
rect 389100 58682 389128 69022
rect 390388 64326 390416 69090
rect 390756 69086 390784 71726
rect 390468 69080 390520 69086
rect 390468 69022 390520 69028
rect 390744 69080 390796 69086
rect 390744 69022 390796 69028
rect 390376 64320 390428 64326
rect 390376 64262 390428 64268
rect 389088 58676 389140 58682
rect 389088 58618 389140 58624
rect 390480 21418 390508 69022
rect 391492 68746 391520 71726
rect 392136 71726 392167 71754
rect 392837 71754 392865 72012
rect 393534 71754 393562 72012
rect 392837 71726 393268 71754
rect 392136 69086 392164 71726
rect 391940 69080 391992 69086
rect 391940 69022 391992 69028
rect 392124 69080 392176 69086
rect 392124 69022 392176 69028
rect 393136 69080 393188 69086
rect 393136 69022 393188 69028
rect 391480 68740 391532 68746
rect 391480 68682 391532 68688
rect 391952 65822 391980 69022
rect 391940 65816 391992 65822
rect 391940 65758 391992 65764
rect 393148 62898 393176 69022
rect 393136 62892 393188 62898
rect 393136 62834 393188 62840
rect 393240 22778 393268 71726
rect 393516 71726 393562 71754
rect 394232 71754 394260 72012
rect 394930 71754 394958 72012
rect 395628 71754 395656 72012
rect 396326 71754 396354 72012
rect 397023 71754 397051 72012
rect 397721 71754 397749 72012
rect 398419 71754 398447 72012
rect 399117 71754 399145 72012
rect 399815 71754 399843 72012
rect 400512 71754 400540 72012
rect 394232 71726 394648 71754
rect 394930 71726 395016 71754
rect 395628 71726 396028 71754
rect 396326 71726 396396 71754
rect 397023 71726 397408 71754
rect 397721 71726 397776 71754
rect 398419 71726 398696 71754
rect 399117 71726 399156 71754
rect 399815 71726 400076 71754
rect 393516 69086 393544 71726
rect 393504 69080 393556 69086
rect 393504 69022 393556 69028
rect 394516 69080 394568 69086
rect 394516 69022 394568 69028
rect 394528 64258 394556 69022
rect 394516 64252 394568 64258
rect 394516 64194 394568 64200
rect 394620 50386 394648 71726
rect 394988 69086 395016 71726
rect 394976 69080 395028 69086
rect 394976 69022 395028 69028
rect 395896 69080 395948 69086
rect 395896 69022 395948 69028
rect 395908 62830 395936 69022
rect 395896 62824 395948 62830
rect 395896 62766 395948 62772
rect 394608 50380 394660 50386
rect 394608 50322 394660 50328
rect 393228 22772 393280 22778
rect 393228 22714 393280 22720
rect 390468 21412 390520 21418
rect 390468 21354 390520 21360
rect 386328 18624 386380 18630
rect 386328 18566 386380 18572
rect 383568 17264 383620 17270
rect 383568 17206 383620 17212
rect 392584 10056 392636 10062
rect 392584 9998 392636 10004
rect 389456 9988 389508 9994
rect 389456 9930 389508 9936
rect 385960 9920 386012 9926
rect 385960 9862 386012 9868
rect 382372 9852 382424 9858
rect 382372 9794 382424 9800
rect 382188 4004 382240 4010
rect 382188 3946 382240 3952
rect 382384 480 382412 9794
rect 384764 8288 384816 8294
rect 384764 8230 384816 8236
rect 383568 3800 383620 3806
rect 383568 3742 383620 3748
rect 383580 480 383608 3742
rect 384776 480 384804 8230
rect 385972 480 386000 9862
rect 388260 8220 388312 8226
rect 388260 8162 388312 8168
rect 387156 3732 387208 3738
rect 387156 3674 387208 3680
rect 387168 480 387196 3674
rect 388272 480 388300 8162
rect 389468 480 389496 9930
rect 391848 8152 391900 8158
rect 391848 8094 391900 8100
rect 390652 3664 390704 3670
rect 390652 3606 390704 3612
rect 390664 480 390692 3606
rect 391860 480 391888 8094
rect 392596 490 392624 9998
rect 395344 8084 395396 8090
rect 395344 8026 395396 8032
rect 394240 3596 394292 3602
rect 394240 3538 394292 3544
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
<<<<<<< HEAD
=======
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 3538
rect 395356 480 395384 8026
rect 396000 3806 396028 71726
rect 396368 69086 396396 71726
rect 396356 69080 396408 69086
rect 396356 69022 396408 69028
rect 397276 69080 397328 69086
rect 397276 69022 397328 69028
rect 396080 10124 396132 10130
rect 396080 10066 396132 10072
rect 395988 3800 396040 3806
rect 395988 3742 396040 3748
rect 396092 490 396120 10066
rect 397288 3874 397316 69022
rect 397380 3942 397408 71726
rect 397748 69086 397776 71726
rect 397736 69080 397788 69086
rect 397736 69022 397788 69028
rect 397368 3936 397420 3942
rect 397368 3878 397420 3884
rect 397276 3868 397328 3874
rect 397276 3810 397328 3816
rect 398668 3670 398696 71726
rect 399128 69086 399156 71726
rect 398748 69080 398800 69086
rect 398748 69022 398800 69028
rect 399116 69080 399168 69086
rect 399116 69022 399168 69028
rect 398760 3738 398788 69022
rect 400048 16574 400076 71726
rect 400508 71726 400540 71754
rect 401210 71754 401238 72012
rect 401908 71754 401936 72012
rect 401210 71726 401456 71754
rect 400508 69086 400536 71726
rect 400128 69080 400180 69086
rect 400128 69022 400180 69028
rect 400496 69080 400548 69086
rect 400496 69022 400548 69028
rect 399956 16546 400076 16574
rect 398840 10192 398892 10198
rect 398840 10134 398892 10140
rect 398748 3732 398800 3738
rect 398748 3674 398800 3680
rect 398656 3664 398708 3670
rect 398656 3606 398708 3612
rect 398852 3534 398880 10134
rect 398932 8016 398984 8022
rect 398932 7958 398984 7964
rect 397736 3528 397788 3534
rect 397736 3470 397788 3476
rect 398840 3528 398892 3534
rect 398840 3470 398892 3476
rect 396368 598 396580 626
rect 396368 490 396396 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 462 396396 490
rect 396552 480 396580 598
rect 397748 480 397776 3470
rect 398944 480 398972 7958
rect 399956 3806 399984 16546
rect 400140 6914 400168 69022
rect 400048 6886 400168 6914
rect 399944 3800 399996 3806
rect 399944 3742 399996 3748
rect 400048 3602 400076 6886
rect 401428 3641 401456 71726
rect 401888 71726 401936 71754
rect 402606 71754 402634 72012
rect 402916 71754 402944 72012
rect 402606 71726 402836 71754
rect 401888 69154 401916 71726
rect 401876 69148 401928 69154
rect 401876 69090 401928 69096
rect 401508 69080 401560 69086
rect 401508 69022 401560 69028
rect 401414 3632 401470 3641
rect 400036 3596 400088 3602
rect 401414 3567 401470 3576
rect 400036 3538 400088 3544
rect 400128 3528 400180 3534
rect 400128 3470 400180 3476
rect 400140 480 400168 3470
rect 401520 3466 401548 69022
rect 402520 7948 402572 7954
rect 402520 7890 402572 7896
rect 401324 3460 401376 3466
rect 401324 3402 401376 3408
rect 401508 3460 401560 3466
rect 401508 3402 401560 3408
rect 401336 480 401364 3402
rect 402532 480 402560 7890
rect 402808 3505 402836 71726
rect 402900 71726 402944 71754
rect 403304 71754 403332 72012
rect 403304 71726 403388 71754
rect 402794 3496 402850 3505
rect 402794 3431 402850 3440
rect 402900 3369 402928 71726
rect 403360 69086 403388 71726
rect 403716 69148 403768 69154
rect 403716 69090 403768 69096
rect 403348 69080 403400 69086
rect 403348 69022 403400 69028
rect 403728 68610 403756 69090
rect 404268 69080 404320 69086
rect 404268 69022 404320 69028
rect 403716 68604 403768 68610
rect 403716 68546 403768 68552
rect 403624 10260 403676 10266
rect 403624 10202 403676 10208
rect 402886 3360 402942 3369
rect 402886 3295 402942 3304
rect 403636 480 403664 10202
rect 404280 3777 404308 69022
rect 406016 7880 406068 7886
rect 406016 7822 406068 7828
rect 404266 3768 404322 3777
rect 404266 3703 404322 3712
rect 404820 2848 404872 2854
rect 404820 2790 404872 2796
rect 404832 480 404860 2790
rect 406028 480 406056 7822
rect 406396 5642 406424 72791
rect 406488 20670 406516 77551
rect 406580 33114 406608 83263
rect 406672 46918 406700 88839
rect 406764 60722 406792 94551
rect 406856 73166 406884 100263
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 406844 73160 406896 73166
rect 406844 73102 406896 73108
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 440240 70372 440292 70378
rect 440240 70314 440292 70320
rect 410524 70100 410576 70106
rect 410524 70042 410576 70048
rect 407120 69420 407172 69426
rect 407120 69362 407172 69368
rect 406752 60716 406804 60722
rect 406752 60658 406804 60664
rect 406660 46912 406712 46918
rect 406660 46854 406712 46860
rect 406568 33108 406620 33114
rect 406568 33050 406620 33056
rect 406476 20664 406528 20670
rect 406476 20606 406528 20612
rect 406384 5636 406436 5642
rect 406384 5578 406436 5584
rect 407132 2922 407160 69362
rect 407212 11008 407264 11014
rect 407212 10950 407264 10956
rect 407120 2916 407172 2922
rect 407120 2858 407172 2864
rect 407224 480 407252 10950
rect 410536 7818 410564 70042
rect 418804 70032 418856 70038
rect 418804 69974 418856 69980
rect 413284 69760 413336 69766
rect 413284 69702 413336 69708
rect 411904 69692 411956 69698
rect 411904 69634 411956 69640
rect 410800 10940 410852 10946
rect 410800 10882 410852 10888
rect 409604 7812 409656 7818
rect 409604 7754 409656 7760
rect 410524 7812 410576 7818
rect 410524 7754 410576 7760
rect 408408 2916 408460 2922
rect 408408 2858 408460 2864
rect 408420 480 408448 2858
rect 409616 480 409644 7754
rect 410812 480 410840 10882
rect 411916 7886 411944 69634
rect 411904 7880 411956 7886
rect 411904 7822 411956 7828
rect 413296 7750 413324 69702
rect 414664 69352 414716 69358
rect 414664 69294 414716 69300
rect 414676 10878 414704 69294
rect 414296 10872 414348 10878
rect 414296 10814 414348 10820
rect 414664 10872 414716 10878
rect 414664 10814 414716 10820
rect 413100 7744 413152 7750
rect 413100 7686 413152 7692
rect 413284 7744 413336 7750
rect 413284 7686 413336 7692
rect 411904 2848 411956 2854
rect 411904 2790 411956 2796
rect 411916 480 411944 2790
rect 413112 480 413140 7686
rect 414308 480 414336 10814
rect 417424 10804 417476 10810
rect 417424 10746 417476 10752
rect 416688 7676 416740 7682
rect 416688 7618 416740 7624
rect 415492 2984 415544 2990
rect 415492 2926 415544 2932
rect 415504 480 415532 2926
rect 416700 480 416728 7618
rect 417436 490 417464 10746
rect 418816 7682 418844 69974
rect 431960 69624 432012 69630
rect 431960 69566 432012 69572
rect 429200 69556 429252 69562
rect 429200 69498 429252 69504
rect 422300 69488 422352 69494
rect 422300 69430 422352 69436
rect 422312 16574 422340 69430
rect 423680 67040 423732 67046
rect 423680 66982 423732 66988
rect 423692 16574 423720 66982
rect 422312 16546 422616 16574
rect 423692 16546 423812 16574
rect 420920 10736 420972 10742
rect 420920 10678 420972 10684
rect 418804 7676 418856 7682
rect 418804 7618 418856 7624
rect 420184 7608 420236 7614
rect 420184 7550 420236 7556
rect 418988 3052 419040 3058
rect 418988 2994 419040 3000
rect 417712 598 417924 626
rect 417712 490 417740 598
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 462 417740 490
rect 417896 480 417924 598
rect 419000 480 419028 2994
rect 420196 480 420224 7550
rect 420932 490 420960 10678
rect 421208 598 421420 626
rect 421208 490 421236 598
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 462 421236 490
rect 421392 480 421420 598
rect 422588 480 422616 16546
rect 423784 480 423812 16546
rect 426808 11960 426860 11966
rect 426808 11902 426860 11908
rect 424968 10668 425020 10674
rect 424968 10610 425020 10616
rect 424980 480 425008 10610
rect 426164 3120 426216 3126
rect 426164 3062 426216 3068
rect 426176 480 426204 3062
rect 426820 490 426848 11902
rect 428464 10600 428516 10606
rect 428464 10542 428516 10548
rect 427096 598 427308 626
rect 427096 490 427124 598
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
<<<<<<< HEAD
rect 427238 -960 427350 480
rect 428434 -960 428546 480
=======
rect 426820 462 427124 490
rect 427280 480 427308 598
rect 428476 480 428504 10542
rect 429212 490 429240 69498
rect 430580 68468 430632 68474
rect 430580 68410 430632 68416
rect 430592 16574 430620 68410
rect 430592 16546 430896 16574
rect 429488 598 429700 626
rect 429488 490 429516 598
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429212 462 429516 490
rect 429672 480 429700 598
rect 430868 480 430896 16546
rect 431972 3126 432000 69566
rect 440252 16574 440280 70314
rect 447140 70304 447192 70310
rect 447140 70246 447192 70252
rect 447152 16574 447180 70246
rect 454040 70236 454092 70242
rect 454040 70178 454092 70184
rect 448520 65612 448572 65618
rect 448520 65554 448572 65560
rect 448532 16574 448560 65554
rect 440252 16546 440372 16574
rect 447152 16546 447456 16574
rect 448532 16546 448652 16574
rect 437480 14476 437532 14482
rect 437480 14418 437532 14424
rect 433984 13252 434036 13258
rect 433984 13194 434036 13200
rect 432052 10532 432104 10538
rect 432052 10474 432104 10480
rect 431960 3120 432012 3126
rect 431960 3062 432012 3068
rect 432064 480 432092 10474
rect 433248 3120 433300 3126
rect 433248 3062 433300 3068
rect 433260 480 433288 3062
rect 433996 490 434024 13194
rect 435088 10464 435140 10470
rect 435088 10406 435140 10412
rect 434272 598 434484 626
rect 434272 490 434300 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 462 434300 490
rect 434456 480 434484 598
rect 435100 490 435128 10406
rect 436744 3188 436796 3194
rect 436744 3130 436796 3136
rect 435376 598 435588 626
rect 435376 490 435404 598
rect 434414 -960 434526 480
rect 435100 462 435404 490
rect 435560 480 435588 598
rect 436756 480 436784 3130
rect 437492 490 437520 14418
rect 439136 10396 439188 10402
rect 439136 10338 439188 10344
rect 437768 598 437980 626
rect 437768 490 437796 598
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437492 462 437796 490
rect 437952 480 437980 598
rect 439148 480 439176 10338
rect 440344 480 440372 16546
rect 441528 15904 441580 15910
rect 441528 15846 441580 15852
rect 441540 480 441568 15846
rect 445760 12164 445812 12170
rect 445760 12106 445812 12112
rect 445024 11824 445076 11830
rect 445024 11766 445076 11772
rect 442632 10328 442684 10334
rect 442632 10270 442684 10276
rect 442644 480 442672 10270
rect 443828 3256 443880 3262
rect 443828 3198 443880 3204
rect 443840 480 443868 3198
rect 445036 480 445064 11766
rect 445772 490 445800 12106
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
<<<<<<< HEAD
=======
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 16546
rect 448624 480 448652 16546
rect 451648 13184 451700 13190
rect 451648 13126 451700 13132
rect 449808 12096 449860 12102
rect 449808 12038 449860 12044
rect 449820 480 449848 12038
rect 450912 3324 450964 3330
rect 450912 3266 450964 3272
rect 450924 480 450952 3266
rect 451660 490 451688 13126
rect 453304 12028 453356 12034
rect 453304 11970 453356 11976
rect 451936 598 452148 626
rect 451936 490 451964 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 462 451964 490
rect 452120 480 452148 598
rect 453316 480 453344 11970
rect 454052 490 454080 70178
rect 460940 70168 460992 70174
rect 460940 70110 460992 70116
rect 456892 64184 456944 64190
rect 456892 64126 456944 64132
rect 455696 9580 455748 9586
rect 455696 9522 455748 9528
rect 454328 598 454540 626
rect 454328 490 454356 598
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 462 454356 490
rect 454512 480 454540 598
rect 455708 480 455736 9522
rect 456904 480 456932 64126
rect 459560 24132 459612 24138
rect 459560 24074 459612 24080
rect 459572 16574 459600 24074
rect 460952 16574 460980 70110
rect 467840 69964 467892 69970
rect 467840 69906 467892 69912
rect 466460 67108 466512 67114
rect 466460 67050 466512 67056
rect 463700 65748 463752 65754
rect 463700 65690 463752 65696
rect 463712 16574 463740 65690
rect 466472 16574 466500 67050
rect 467852 16574 467880 69906
rect 474740 69896 474792 69902
rect 474740 69838 474792 69844
rect 472624 69828 472676 69834
rect 472624 69770 472676 69776
rect 470600 65680 470652 65686
rect 470600 65622 470652 65628
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 463712 16546 464016 16574
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 459192 9444 459244 9450
rect 459192 9386 459244 9392
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 9386
rect 459940 490 459968 16546
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
<<<<<<< HEAD
=======
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 16546
rect 462780 9376 462832 9382
rect 462780 9318 462832 9324
rect 462792 480 462820 9318
rect 463988 480 464016 16546
rect 466276 9172 466328 9178
rect 466276 9114 466328 9120
rect 465172 4140 465224 4146
rect 465172 4082 465224 4088
rect 465184 480 465212 4082
rect 466288 480 466316 9114
rect 467484 480 467512 16546
rect 468220 490 468248 16546
rect 469864 9104 469916 9110
rect 469864 9046 469916 9052
rect 468496 598 468708 626
rect 468496 490 468524 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 462 468524 490
rect 468680 480 468708 598
rect 469876 480 469904 9046
rect 470612 490 470640 65622
rect 472636 4214 472664 69770
rect 474752 16574 474780 69838
rect 492680 68876 492732 68882
rect 492680 68818 492732 68824
rect 481640 68672 481692 68678
rect 481640 68614 481692 68620
rect 474752 16546 475792 16574
rect 473452 9036 473504 9042
rect 473452 8978 473504 8984
rect 472624 4208 472676 4214
rect 472624 4150 472676 4156
rect 472256 4072 472308 4078
rect 472256 4014 472308 4020
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 468638 -960 468750 480
rect 469834 -960 469946 480
<<<<<<< HEAD
=======
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 4014
rect 473464 480 473492 8978
rect 474556 4208 474608 4214
rect 474556 4150 474608 4156
rect 474568 480 474596 4150
rect 475764 480 475792 16546
rect 478144 14544 478196 14550
rect 478144 14486 478196 14492
rect 476948 8968 477000 8974
rect 476948 8910 477000 8916
rect 476960 480 476988 8910
rect 478156 480 478184 14486
rect 480536 7880 480588 7886
rect 480536 7822 480588 7828
rect 479340 4004 479392 4010
rect 479340 3946 479392 3952
rect 479352 480 479380 3946
rect 480548 480 480576 7822
rect 481652 6914 481680 68614
rect 488540 68536 488592 68542
rect 488540 68478 488592 68484
rect 483020 68400 483072 68406
rect 483020 68342 483072 68348
rect 481732 17264 481784 17270
rect 481732 17206 481784 17212
rect 481744 16574 481772 17206
rect 483032 16574 483060 68342
rect 484400 67176 484452 67182
rect 484400 67118 484452 67124
rect 484412 16574 484440 67118
rect 485780 64388 485832 64394
rect 485780 64330 485832 64336
rect 485792 16574 485820 64330
rect 488552 16574 488580 68478
rect 489920 66972 489972 66978
rect 489920 66914 489972 66920
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 482388 490 482416 16546
rect 482664 598 482876 626
rect 482664 490 482692 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
<<<<<<< HEAD
=======
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 16546
rect 484780 490 484808 16546
rect 485056 598 485268 626
rect 485056 490 485084 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 462 485084 490
rect 485240 480 485268 598
rect 486436 480 486464 16546
rect 487620 7336 487672 7342
rect 487620 7278 487672 7284
rect 487632 480 487660 7278
rect 488828 480 488856 16546
rect 489932 4010 489960 66914
rect 492692 16574 492720 68818
rect 503720 68808 503772 68814
rect 503720 68750 503772 68756
rect 500960 68332 501012 68338
rect 500960 68274 501012 68280
rect 496820 67312 496872 67318
rect 496820 67254 496872 67260
rect 496832 16574 496860 67254
rect 499580 18624 499632 18630
rect 499580 18566 499632 18572
rect 499592 16574 499620 18566
rect 500972 16574 501000 68274
rect 492692 16546 493088 16574
rect 496832 16546 497136 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 490012 10872 490064 10878
rect 490012 10814 490064 10820
rect 489920 4004 489972 4010
rect 489920 3946 489972 3952
rect 490024 3482 490052 10814
rect 492312 7676 492364 7682
rect 492312 7618 492364 7624
rect 491116 4004 491168 4010
rect 491116 3946 491168 3952
rect 489932 3454 490052 3482
rect 489932 480 489960 3454
rect 491128 480 491156 3946
rect 492324 480 492352 7618
rect 493060 490 493088 16546
rect 494704 13116 494756 13122
rect 494704 13058 494756 13064
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
<<<<<<< HEAD
=======
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 13058
rect 495900 7812 495952 7818
rect 495900 7754 495952 7760
rect 495912 480 495940 7754
rect 497108 480 497136 16546
rect 498936 11892 498988 11898
rect 498936 11834 498988 11840
rect 498200 11756 498252 11762
rect 498200 11698 498252 11704
rect 498212 480 498240 11698
rect 498948 490 498976 11834
rect 499224 598 499436 626
rect 499224 490 499252 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 462 499252 490
rect 499408 480 499436 598
rect 500604 480 500632 16546
rect 501340 490 501368 16546
rect 502984 5704 503036 5710
rect 502984 5646 503036 5652
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 499366 -960 499478 480
rect 500562 -960 500674 480
<<<<<<< HEAD
=======
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 5646
rect 503732 490 503760 68750
rect 528560 68740 528612 68746
rect 528560 68682 528612 68688
rect 506480 67244 506532 67250
rect 506480 67186 506532 67192
rect 506492 16574 506520 67186
rect 507860 66904 507912 66910
rect 507860 66846 507912 66852
rect 507872 16574 507900 66846
rect 510620 65884 510672 65890
rect 510620 65826 510672 65832
rect 510632 16574 510660 65826
rect 524420 65816 524472 65822
rect 524420 65758 524472 65764
rect 517520 64320 517572 64326
rect 517520 64262 517572 64268
rect 514760 58676 514812 58682
rect 514760 58618 514812 58624
rect 506492 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 505376 7744 505428 7750
rect 505376 7686 505428 7692
rect 504008 598 504220 626
rect 504008 490 504036 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 462 504036 490
rect 504192 480 504220 598
rect 505388 480 505416 7686
rect 506480 5772 506532 5778
rect 506480 5714 506532 5720
rect 506492 480 506520 5714
rect 507228 490 507256 16546
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
<<<<<<< HEAD
=======
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 16546
rect 510068 5840 510120 5846
rect 510068 5782 510120 5788
rect 510080 480 510108 5782
rect 511276 480 511304 16546
rect 513564 5908 513616 5914
rect 513564 5850 513616 5856
rect 512460 4344 512512 4350
rect 512460 4286 512512 4292
rect 512472 480 512500 4286
rect 513576 480 513604 5850
rect 514772 480 514800 58618
rect 517532 16574 517560 64262
rect 521660 21412 521712 21418
rect 521660 21354 521712 21360
rect 521672 16574 521700 21354
rect 524432 16574 524460 65758
rect 517532 16546 517928 16574
rect 521672 16546 521884 16574
rect 524432 16546 525472 16574
rect 517152 5976 517204 5982
rect 517152 5918 517204 5924
rect 515956 4412 516008 4418
rect 515956 4354 516008 4360
rect 515968 480 515996 4354
rect 517164 480 517192 5918
rect 517900 490 517928 16546
rect 520740 6044 520792 6050
rect 520740 5986 520792 5992
rect 519544 4480 519596 4486
rect 519544 4422 519596 4428
rect 518176 598 518388 626
rect 518176 490 518204 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
<<<<<<< HEAD
=======
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 4422
rect 520752 480 520780 5986
rect 521856 480 521884 16546
rect 524236 6112 524288 6118
rect 524236 6054 524288 6060
rect 523040 4548 523092 4554
rect 523040 4490 523092 4496
rect 523052 480 523080 4490
rect 524248 480 524276 6054
rect 525444 480 525472 16546
rect 527824 6860 527876 6866
rect 527824 6802 527876 6808
rect 526628 4616 526680 4622
rect 526628 4558 526680 4564
rect 526640 480 526668 4558
rect 527836 480 527864 6802
rect 528572 490 528600 68682
rect 579620 68604 579672 68610
rect 579620 68546 579672 68552
rect 575480 65544 575532 65550
rect 575480 65486 575532 65492
rect 539600 64252 539652 64258
rect 539600 64194 539652 64200
rect 530584 62892 530636 62898
rect 530584 62834 530636 62840
rect 530124 4684 530176 4690
rect 530124 4626 530176 4632
rect 528848 598 529060 626
rect 528848 490 528876 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
<<<<<<< HEAD
=======
rect 528572 462 528876 490
rect 529032 480 529060 598
rect 530136 480 530164 4626
rect 530596 3398 530624 62834
rect 535460 22772 535512 22778
rect 535460 22714 535512 22720
rect 535472 16574 535500 22714
rect 535472 16546 536144 16574
rect 531320 6792 531372 6798
rect 531320 6734 531372 6740
rect 530584 3392 530636 3398
rect 530584 3334 530636 3340
rect 531332 480 531360 6734
rect 534908 6724 534960 6730
rect 534908 6666 534960 6672
rect 533712 4752 533764 4758
rect 533712 4694 533764 4700
rect 532516 3392 532568 3398
rect 532516 3334 532568 3340
rect 532528 480 532556 3334
rect 533724 480 533752 4694
rect 534920 480 534948 6666
rect 536116 480 536144 16546
rect 538404 6656 538456 6662
rect 538404 6598 538456 6604
rect 537208 5500 537260 5506
rect 537208 5442 537260 5448
rect 537220 480 537248 5442
rect 538416 480 538444 6598
rect 539612 480 539640 64194
rect 546500 62824 546552 62830
rect 546500 62766 546552 62772
rect 542360 50380 542412 50386
rect 542360 50322 542412 50328
rect 542372 16574 542400 50322
rect 546512 16574 546540 62766
rect 575492 16574 575520 65486
rect 579632 16574 579660 68546
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 579894 33144 579950 33153
rect 579894 33079 579896 33088
rect 579948 33079 579950 33088
rect 579896 33050 579948 33056
rect 579896 20664 579948 20670
rect 579896 20606 579948 20612
rect 579908 19825 579936 20606
rect 579894 19816 579950 19825
rect 579894 19751 579950 19760
rect 542372 16546 542768 16574
rect 546512 16546 546724 16574
rect 575492 16546 575888 16574
rect 579632 16546 579844 16574
rect 541992 6588 542044 6594
rect 541992 6530 542044 6536
rect 540796 5432 540848 5438
rect 540796 5374 540848 5380
rect 540808 480 540836 5374
rect 542004 480 542032 6530
rect 542740 490 542768 16546
rect 545488 6520 545540 6526
rect 545488 6462 545540 6468
rect 544384 5364 544436 5370
rect 544384 5306 544436 5312
rect 543016 598 543228 626
rect 543016 490 543044 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
<<<<<<< HEAD
=======
rect 542740 462 543044 490
rect 543200 480 543228 598
rect 544396 480 544424 5306
rect 545500 480 545528 6462
rect 546696 480 546724 16546
rect 563244 9648 563296 9654
rect 563244 9590 563296 9596
rect 549076 6452 549128 6458
rect 549076 6394 549128 6400
rect 547880 5296 547932 5302
rect 547880 5238 547932 5244
rect 547892 480 547920 5238
rect 549088 480 549116 6394
rect 552664 6384 552716 6390
rect 552664 6326 552716 6332
rect 551468 5228 551520 5234
rect 551468 5170 551520 5176
rect 550272 3936 550324 3942
rect 550272 3878 550324 3884
rect 550284 480 550312 3878
rect 551480 480 551508 5170
rect 552676 480 552704 6326
rect 556160 6316 556212 6322
rect 556160 6258 556212 6264
rect 554964 5160 555016 5166
rect 554964 5102 555016 5108
rect 553768 3868 553820 3874
rect 553768 3810 553820 3816
rect 553780 480 553808 3810
rect 554976 480 555004 5102
rect 556172 480 556200 6258
rect 559748 6248 559800 6254
rect 559748 6190 559800 6196
rect 558552 5092 558604 5098
rect 558552 5034 558604 5040
rect 557356 3800 557408 3806
rect 557356 3742 557408 3748
rect 557368 480 557396 3742
rect 558564 480 558592 5034
rect 559760 480 559788 6190
rect 562048 5024 562100 5030
rect 562048 4966 562100 4972
rect 560852 3732 560904 3738
rect 560852 3674 560904 3680
rect 560864 480 560892 3674
rect 562060 480 562088 4966
rect 563256 480 563284 9590
rect 570328 9512 570380 9518
rect 570328 9454 570380 9460
rect 566832 6180 566884 6186
rect 566832 6122 566884 6128
rect 565636 4956 565688 4962
rect 565636 4898 565688 4904
rect 564440 3664 564492 3670
rect 564440 3606 564492 3612
rect 564452 480 564480 3606
rect 565648 480 565676 4898
rect 566844 480 566872 6122
rect 569132 4888 569184 4894
rect 569132 4830 569184 4836
rect 568028 3596 568080 3602
rect 568028 3538 568080 3544
rect 568040 480 568068 3538
rect 569144 480 569172 4830
rect 570340 480 570368 9454
rect 573916 9308 573968 9314
rect 573916 9250 573968 9256
rect 572720 4820 572772 4826
rect 572720 4762 572772 4768
rect 571524 3528 571576 3534
rect 571524 3470 571576 3476
rect 571536 480 571564 3470
rect 572732 480 572760 4762
rect 573928 480 573956 9250
rect 575112 3460 575164 3466
rect 575112 3402 575164 3408
rect 575124 480 575152 3402
rect 575860 490 575888 16546
rect 577412 9240 577464 9246
rect 577412 9182 577464 9188
rect 576136 598 576348 626
rect 576136 490 576164 598
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 462 576164 490
rect 576320 480 576348 598
rect 577424 480 577452 9182
rect 578606 3632 578662 3641
rect 578606 3567 578662 3576
rect 578620 480 578648 3567
rect 579816 480 579844 16546
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 580184 5642 580212 6559
rect 580172 5636 580224 5642
rect 580172 5578 580224 5584
rect 582194 3768 582250 3777
rect 582194 3703 582250 3712
rect 580998 3496 581054 3505
rect 580998 3431 581054 3440
rect 581012 480 581040 3431
rect 582208 480 582236 3703
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 697312 3478 697368
rect 3146 684256 3202 684312
rect 3146 658144 3202 658200
rect 3330 632068 3332 632088
rect 3332 632068 3384 632088
rect 3384 632068 3386 632088
rect 3330 632032 3386 632068
rect 2962 619112 3018 619168
rect 3330 606056 3386 606112
rect 2778 593000 2834 593056
rect 3330 579944 3386 580000
rect 3054 566888 3110 566944
rect 3330 553832 3386 553888
rect 3330 540776 3386 540832
rect 3330 527856 3386 527912
rect 3238 501744 3294 501800
rect 2870 475632 2926 475688
rect 3054 462576 3110 462632
rect 2962 449520 3018 449576
rect 2962 423544 3018 423600
rect 3330 384376 3386 384432
rect 3238 371320 3294 371376
rect 3146 319232 3202 319288
rect 3054 306176 3110 306232
rect 2962 293120 3018 293176
rect 2870 254088 2926 254144
rect 3514 671200 3570 671256
rect 3422 358400 3478 358456
rect 3606 645088 3662 645144
rect 3514 345344 3570 345400
rect 3698 514800 3754 514856
rect 3606 332288 3662 332344
rect 3422 214920 3478 214976
rect 3790 488688 3846 488744
rect 3698 280064 3754 280120
rect 3514 201864 3570 201920
rect 3882 436600 3938 436656
rect 3790 267144 3846 267200
rect 3606 188808 3662 188864
rect 3974 410488 4030 410544
rect 4066 397432 4122 397488
rect 3882 241032 3938 241088
rect 3698 175888 3754 175944
rect 3422 149776 3478 149832
rect 580170 697176 580226 697232
rect 57426 365064 57482 365120
rect 406014 364964 406016 364984
rect 406016 364964 406068 364984
rect 406068 364964 406070 364984
rect 406014 364928 406070 364964
rect 57150 360440 57206 360496
rect 57242 354864 57298 354920
rect 57610 349288 57666 349344
rect 57610 343712 57666 343768
rect 57610 338272 57666 338328
rect 57610 332696 57666 332752
rect 57334 327120 57390 327176
rect 57334 321544 57390 321600
rect 57610 316104 57666 316160
rect 57610 310428 57612 310448
rect 57612 310428 57664 310448
rect 57664 310428 57666 310448
rect 57610 310392 57666 310428
rect 57426 304972 57482 305008
rect 57426 304952 57428 304972
rect 57428 304952 57480 304972
rect 57480 304952 57482 304972
rect 57610 299412 57612 299432
rect 57612 299412 57664 299432
rect 57664 299412 57666 299432
rect 57610 299376 57666 299412
rect 405830 298152 405886 298208
rect 57610 293800 57666 293856
rect 57610 288380 57666 288416
rect 57610 288360 57612 288380
rect 57612 288360 57664 288380
rect 57664 288360 57666 288380
rect 57610 282820 57612 282840
rect 57612 282820 57664 282840
rect 57664 282820 57666 282840
rect 57610 282784 57666 282820
rect 57610 277208 57666 277264
rect 57518 271632 57574 271688
rect 57334 266056 57390 266112
rect 57426 260616 57482 260672
rect 57610 255040 57666 255096
rect 57242 249464 57298 249520
rect 57426 243888 57482 243944
rect 57610 238448 57666 238504
rect 57610 232872 57666 232928
rect 406382 360304 406438 360360
rect 406474 354592 406530 354648
rect 406290 247152 406346 247208
rect 406198 241576 406254 241632
rect 406106 230288 406162 230344
rect 3974 227976 4030 228032
rect 57610 227296 57666 227352
rect 406290 224612 406292 224632
rect 406292 224612 406344 224632
rect 406344 224612 406346 224632
rect 406290 224576 406346 224612
rect 57610 221720 57666 221776
rect 406474 349052 406476 349072
rect 406476 349052 406528 349072
rect 406528 349052 406530 349072
rect 406474 349016 406530 349052
rect 406474 343340 406476 343360
rect 406476 343340 406528 343360
rect 406528 343340 406530 343360
rect 406474 343304 406530 343340
rect 406474 337728 406530 337784
rect 406474 332016 406530 332072
rect 406566 326304 406622 326360
rect 406382 219000 406438 219056
rect 57058 216144 57114 216200
rect 56782 210704 56838 210760
rect 57610 205128 57666 205184
rect 57610 199552 57666 199608
rect 57610 193976 57666 194032
rect 57610 188536 57666 188592
rect 57610 182960 57666 183016
rect 56690 177384 56746 177440
rect 57610 171808 57666 171864
rect 57610 166232 57666 166288
rect 3790 162832 3846 162888
rect 406382 213288 406438 213344
rect 406658 320728 406714 320784
rect 406750 315016 406806 315072
rect 406474 207712 406530 207768
rect 406290 162424 406346 162480
rect 57610 160792 57666 160848
rect 406842 309440 406898 309496
rect 406842 303728 406898 303784
rect 406566 202000 406622 202056
rect 406842 292476 406844 292496
rect 406844 292476 406896 292496
rect 406896 292476 406898 292496
rect 406842 292440 406898 292476
rect 406842 286728 406898 286784
rect 406842 281152 406898 281208
rect 406934 275440 406990 275496
rect 406658 196288 406714 196344
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580262 657328 580318 657384
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 407026 269864 407082 269920
rect 407026 264152 407082 264208
rect 406382 156712 406438 156768
rect 57610 155216 57666 155272
rect 56874 149640 56930 149696
rect 57518 144064 57574 144120
rect 57518 138488 57574 138544
rect 3514 136720 3570 136776
rect 406750 190712 406806 190768
rect 406658 185000 406714 185056
rect 406934 258032 406990 258088
rect 407026 252884 407082 252920
rect 407026 252864 407028 252884
rect 407028 252864 407080 252884
rect 407080 252864 407082 252884
rect 406842 179424 406898 179480
rect 406474 151136 406530 151192
rect 407026 235900 407028 235920
rect 407028 235900 407080 235920
rect 407080 235900 407082 235920
rect 407026 235864 407082 235900
rect 406934 173712 406990 173768
rect 580170 617480 580226 617536
rect 579618 590960 579674 591016
rect 579618 577632 579674 577688
rect 579894 564304 579950 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 579618 484608 579674 484664
rect 579986 471416 580042 471472
rect 579986 431568 580042 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 579802 378392 579858 378448
rect 580170 365064 580226 365120
rect 580354 604152 580410 604208
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580262 338544 580318 338600
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245520 580226 245576
rect 579618 232328 579674 232384
rect 580170 219000 580226 219056
rect 580446 551112 580502 551168
rect 580538 511264 580594 511320
rect 580630 497936 580686 497992
rect 580354 285368 580410 285424
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 580170 192480 580226 192536
rect 580722 458088 580778 458144
rect 580814 444760 580870 444816
rect 580906 391720 580962 391776
rect 580170 179152 580226 179208
rect 407026 168136 407082 168192
rect 580170 165824 580226 165880
rect 406566 145424 406622 145480
rect 579986 152632 580042 152688
rect 406658 139848 406714 139904
rect 580170 139304 580226 139360
rect 406382 134136 406438 134192
rect 57518 133048 57574 133104
rect 406474 128560 406530 128616
rect 56966 127472 57022 127528
rect 580170 125976 580226 126032
rect 3606 123664 3662 123720
rect 407026 122848 407082 122904
rect 57058 121896 57114 121952
rect 406382 117136 406438 117192
rect 57610 116320 57666 116376
rect 579802 112784 579858 112840
rect 406474 111560 406530 111616
rect 57610 110744 57666 110800
rect 3422 110608 3478 110664
rect 406382 105848 406438 105904
rect 57426 105168 57482 105224
rect 57426 99728 57482 99784
rect 3514 97552 3570 97608
rect 3422 84632 3478 84688
rect 57610 94152 57666 94208
rect 57518 88576 57574 88632
rect 406842 100272 406898 100328
rect 406750 94560 406806 94616
rect 406658 88848 406714 88904
rect 406566 83272 406622 83328
rect 57426 83000 57482 83056
rect 57518 77560 57574 77616
rect 406474 77560 406530 77616
rect 57426 72800 57482 72856
rect 406382 72800 406438 72856
rect 3882 71576 3938 71632
rect 3790 58520 3846 58576
rect 3698 45464 3754 45520
rect 3606 32408 3662 32464
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 5262 3304 5318 3360
rect 11150 3440 11206 3496
rect 20626 3576 20682 3632
rect 25318 3712 25374 3768
rect 131210 3712 131266 3768
rect 131118 3576 131174 3632
rect 129830 3440 129886 3496
rect 132590 3304 132646 3360
rect 138846 3304 138902 3360
rect 142434 3440 142490 3496
rect 241702 3576 241758 3632
rect 245198 3712 245254 3768
rect 314750 3440 314806 3496
rect 314842 3304 314898 3360
rect 333978 3576 334034 3632
rect 335542 3712 335598 3768
rect 401414 3576 401470 3632
rect 402794 3440 402850 3496
rect 402886 3304 402942 3360
rect 404266 3712 404322 3768
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 579894 33108 579950 33144
rect 579894 33088 579896 33108
rect 579896 33088 579948 33108
rect 579948 33088 579950 33108
rect 579894 19760 579950 19816
rect 578606 3576 578662 3632
rect 580170 6568 580226 6624
rect 582194 3712 582250 3768
rect 580998 3440 581054 3496
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697370 480 697460
rect 3417 697370 3483 697373
rect -960 697368 3483 697370
rect -960 697312 3422 697368
rect 3478 697312 3483 697368
rect -960 697310 3483 697312
rect -960 697220 480 697310
rect 3417 697307 3483 697310
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3141 684314 3207 684317
rect -960 684312 3207 684314
rect -960 684256 3146 684312
rect 3202 684256 3207 684312
rect -960 684254 3207 684256
rect -960 684164 480 684254
rect 3141 684251 3207 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3141 658202 3207 658205
rect -960 658200 3207 658202
rect -960 658144 3146 658200
rect 3202 658144 3207 658200
rect -960 658142 3207 658144
rect -960 658052 480 658142
rect 3141 658139 3207 658142
rect 580257 657386 580323 657389
rect 583520 657386 584960 657476
rect 580257 657384 584960 657386
rect 580257 657328 580262 657384
rect 580318 657328 584960 657384
rect 580257 657326 584960 657328
rect 580257 657323 580323 657326
rect 583520 657236 584960 657326
rect -960 645146 480 645236
rect 3601 645146 3667 645149
rect -960 645144 3667 645146
rect -960 645088 3606 645144
rect 3662 645088 3667 645144
rect -960 645086 3667 645088
rect -960 644996 480 645086
rect 3601 645083 3667 645086
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3325 632090 3391 632093
rect -960 632088 3391 632090
rect -960 632032 3330 632088
rect 3386 632032 3391 632088
rect -960 632030 3391 632032
rect -960 631940 480 632030
rect 3325 632027 3391 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 2957 619170 3023 619173
rect -960 619168 3023 619170
rect -960 619112 2962 619168
rect 3018 619112 3023 619168
rect -960 619110 3023 619112
rect -960 619020 480 619110
rect 2957 619107 3023 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 580349 604210 580415 604213
rect 583520 604210 584960 604300
rect 580349 604208 584960 604210
rect 580349 604152 580354 604208
rect 580410 604152 584960 604208
rect 580349 604150 584960 604152
rect 580349 604147 580415 604150
rect 583520 604060 584960 604150
rect -960 593058 480 593148
rect 2773 593058 2839 593061
rect -960 593056 2839 593058
rect -960 593000 2778 593056
rect 2834 593000 2839 593056
rect -960 592998 2839 593000
rect -960 592908 480 592998
rect 2773 592995 2839 592998
rect 579613 591018 579679 591021
rect 583520 591018 584960 591108
rect 579613 591016 584960 591018
rect 579613 590960 579618 591016
rect 579674 590960 584960 591016
rect 579613 590958 584960 590960
rect 579613 590955 579679 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 579889 564362 579955 564365
rect 583520 564362 584960 564452
rect 579889 564360 584960 564362
rect 579889 564304 579894 564360
rect 579950 564304 584960 564360
rect 579889 564302 584960 564304
rect 579889 564299 579955 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 580441 551170 580507 551173
rect 583520 551170 584960 551260
rect 580441 551168 584960 551170
rect 580441 551112 580446 551168
rect 580502 551112 584960 551168
rect 580441 551110 584960 551112
rect 580441 551107 580507 551110
rect 583520 551020 584960 551110
rect -960 540834 480 540924
rect 3325 540834 3391 540837
rect -960 540832 3391 540834
rect -960 540776 3330 540832
rect 3386 540776 3391 540832
rect -960 540774 3391 540776
rect -960 540684 480 540774
rect 3325 540771 3391 540774
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3693 514858 3759 514861
rect -960 514856 3759 514858
rect -960 514800 3698 514856
rect 3754 514800 3759 514856
rect -960 514798 3759 514800
rect -960 514708 480 514798
rect 3693 514795 3759 514798
rect 580533 511322 580599 511325
rect 583520 511322 584960 511412
rect 580533 511320 584960 511322
rect 580533 511264 580538 511320
rect 580594 511264 584960 511320
rect 580533 511262 584960 511264
rect 580533 511259 580599 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 580625 497994 580691 497997
rect 583520 497994 584960 498084
rect 580625 497992 584960 497994
rect 580625 497936 580630 497992
rect 580686 497936 584960 497992
rect 580625 497934 584960 497936
rect 580625 497931 580691 497934
rect 583520 497844 584960 497934
rect -960 488746 480 488836
rect 3785 488746 3851 488749
rect -960 488744 3851 488746
rect -960 488688 3790 488744
rect 3846 488688 3851 488744
rect -960 488686 3851 488688
rect -960 488596 480 488686
rect 3785 488683 3851 488686
rect 579613 484666 579679 484669
rect 583520 484666 584960 484756
rect 579613 484664 584960 484666
rect 579613 484608 579618 484664
rect 579674 484608 584960 484664
rect 579613 484606 584960 484608
rect 579613 484603 579679 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 2865 475690 2931 475693
rect -960 475688 2931 475690
rect -960 475632 2870 475688
rect 2926 475632 2931 475688
rect -960 475630 2931 475632
rect -960 475540 480 475630
rect 2865 475627 2931 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3049 462634 3115 462637
rect -960 462632 3115 462634
rect -960 462576 3054 462632
rect 3110 462576 3115 462632
rect -960 462574 3115 462576
rect -960 462484 480 462574
rect 3049 462571 3115 462574
rect 580717 458146 580783 458149
rect 583520 458146 584960 458236
rect 580717 458144 584960 458146
rect 580717 458088 580722 458144
rect 580778 458088 584960 458144
rect 580717 458086 584960 458088
rect 580717 458083 580783 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 2957 449578 3023 449581
rect -960 449576 3023 449578
rect -960 449520 2962 449576
rect 3018 449520 3023 449576
rect -960 449518 3023 449520
rect -960 449428 480 449518
rect 2957 449515 3023 449518
rect 580809 444818 580875 444821
rect 583520 444818 584960 444908
rect 580809 444816 584960 444818
rect 580809 444760 580814 444816
rect 580870 444760 584960 444816
rect 580809 444758 584960 444760
rect 580809 444755 580875 444758
rect 583520 444668 584960 444758
rect -960 436658 480 436748
rect 3877 436658 3943 436661
rect -960 436656 3943 436658
rect -960 436600 3882 436656
rect 3938 436600 3943 436656
rect -960 436598 3943 436600
rect -960 436508 480 436598
rect 3877 436595 3943 436598
rect 579981 431626 580047 431629
rect 583520 431626 584960 431716
rect 579981 431624 584960 431626
rect 579981 431568 579986 431624
rect 580042 431568 584960 431624
rect 579981 431566 584960 431568
rect 579981 431563 580047 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2957 423602 3023 423605
rect -960 423600 3023 423602
rect -960 423544 2962 423600
rect 3018 423544 3023 423600
rect -960 423542 3023 423544
rect -960 423452 480 423542
rect 2957 423539 3023 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3969 410546 4035 410549
rect -960 410544 4035 410546
rect -960 410488 3974 410544
rect 4030 410488 4035 410544
rect -960 410486 4035 410488
rect -960 410396 480 410486
rect 3969 410483 4035 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 4061 397490 4127 397493
rect -960 397488 4127 397490
rect -960 397432 4066 397488
rect 4122 397432 4127 397488
rect -960 397430 4127 397432
rect -960 397340 480 397430
rect 4061 397427 4127 397430
rect 580901 391778 580967 391781
rect 583520 391778 584960 391868
rect 580901 391776 584960 391778
rect 580901 391720 580906 391776
rect 580962 391720 584960 391776
rect 580901 391718 584960 391720
rect 580901 391715 580967 391718
rect 583520 391628 584960 391718
rect -960 384434 480 384524
rect 3325 384434 3391 384437
rect -960 384432 3391 384434
rect -960 384376 3330 384432
rect 3386 384376 3391 384432
rect -960 384374 3391 384376
rect -960 384284 480 384374
rect 3325 384371 3391 384374
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 579797 378387 579863 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect -960 371318 3299 371320
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 57421 365122 57487 365125
rect 59494 365122 60076 365128
rect 57421 365120 60076 365122
rect 57421 365064 57426 365120
rect 57482 365068 60076 365120
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 57482 365064 59554 365068
rect 57421 365062 59554 365064
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 57421 365059 57487 365062
rect 580165 365059 580231 365062
rect 404064 364986 404738 365006
rect 406009 364986 406075 364989
rect 404064 364984 406075 364986
rect 404064 364946 406014 364984
rect 404678 364928 406014 364946
rect 406070 364928 406075 364984
rect 583520 364972 584960 365062
rect 404678 364926 406075 364928
rect 406009 364923 406075 364926
rect 57145 360498 57211 360501
rect 57145 360496 59554 360498
rect 57145 360440 57150 360496
rect 57206 360443 59554 360496
rect 57206 360440 60076 360443
rect 57145 360438 60076 360440
rect 57145 360435 57211 360438
rect 59494 360383 60076 360438
rect 406377 360362 406443 360365
rect 404678 360360 406443 360362
rect 404678 360333 406382 360360
rect 404064 360304 406382 360333
rect 406438 360304 406443 360360
rect 404064 360302 406443 360304
rect 404064 360273 404738 360302
rect 406377 360299 406443 360302
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 57237 354922 57303 354925
rect 57237 354920 59554 354922
rect 57237 354864 57242 354920
rect 57298 354896 59554 354920
rect 57298 354864 60076 354896
rect 57237 354862 60076 354864
rect 57237 354859 57303 354862
rect 59494 354836 60076 354862
rect 404064 354650 404738 354680
rect 406469 354650 406535 354653
rect 404064 354648 406535 354650
rect 404064 354620 406474 354648
rect 404678 354592 406474 354620
rect 406530 354592 406535 354648
rect 404678 354590 406535 354592
rect 406469 354587 406535 354590
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 57605 349346 57671 349349
rect 59494 349346 60076 349350
rect 57605 349344 60076 349346
rect 57605 349288 57610 349344
rect 57666 349290 60076 349344
rect 57666 349288 59554 349290
rect 57605 349286 59554 349288
rect 57605 349283 57671 349286
rect 406469 349074 406535 349077
rect 404678 349072 406535 349074
rect 404678 349027 406474 349072
rect 404064 349016 406474 349027
rect 406530 349016 406535 349072
rect 404064 349014 406535 349016
rect 404064 348967 404738 349014
rect 406469 349011 406535 349014
rect -960 345402 480 345492
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 57605 343770 57671 343773
rect 59494 343770 60076 343804
rect 57605 343768 60076 343770
rect 57605 343712 57610 343768
rect 57666 343744 60076 343768
rect 57666 343712 59554 343744
rect 57605 343710 59554 343712
rect 57605 343707 57671 343710
rect 404064 343362 404738 343374
rect 406469 343362 406535 343365
rect 404064 343360 406535 343362
rect 404064 343314 406474 343360
rect 404678 343304 406474 343314
rect 406530 343304 406535 343360
rect 404678 343302 406535 343304
rect 406469 343299 406535 343302
rect 580257 338602 580323 338605
rect 583520 338602 584960 338692
rect 580257 338600 584960 338602
rect 580257 338544 580262 338600
rect 580318 338544 584960 338600
rect 580257 338542 584960 338544
rect 580257 338539 580323 338542
rect 583520 338452 584960 338542
rect 57605 338330 57671 338333
rect 57605 338328 59554 338330
rect 57605 338272 57610 338328
rect 57666 338272 59554 338328
rect 57605 338270 59554 338272
rect 57605 338267 57671 338270
rect 59494 338257 59554 338270
rect 59494 338197 60076 338257
rect 406469 337786 406535 337789
rect 404310 337784 406535 337786
rect 404310 337728 406474 337784
rect 406530 337728 406535 337784
rect 404310 337726 406535 337728
rect 404310 337721 404370 337726
rect 406469 337723 406535 337726
rect 404064 337661 404370 337721
rect 57605 332754 57671 332757
rect 57605 332752 59554 332754
rect 57605 332696 57610 332752
rect 57666 332711 59554 332752
rect 57666 332696 60076 332711
rect 57605 332694 60076 332696
rect 57605 332691 57671 332694
rect 59494 332651 60076 332694
rect -960 332346 480 332436
rect 3601 332346 3667 332349
rect -960 332344 3667 332346
rect -960 332288 3606 332344
rect 3662 332288 3667 332344
rect -960 332286 3667 332288
rect -960 332196 480 332286
rect 3601 332283 3667 332286
rect 406469 332074 406535 332077
rect 404678 332072 406535 332074
rect 404678 332068 406474 332072
rect 404064 332016 406474 332068
rect 406530 332016 406535 332072
rect 404064 332014 406535 332016
rect 404064 332008 404738 332014
rect 406469 332011 406535 332014
rect 57329 327178 57395 327181
rect 57329 327176 59554 327178
rect 57329 327120 57334 327176
rect 57390 327164 59554 327176
rect 57390 327120 60076 327164
rect 57329 327118 60076 327120
rect 57329 327115 57395 327118
rect 59494 327104 60076 327118
rect 404064 326362 404738 326415
rect 406561 326362 406627 326365
rect 404064 326360 406627 326362
rect 404064 326355 406566 326360
rect 404678 326304 406566 326355
rect 406622 326304 406627 326360
rect 404678 326302 406627 326304
rect 406561 326299 406627 326302
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 57329 321602 57395 321605
rect 59494 321602 60076 321618
rect 57329 321600 60076 321602
rect 57329 321544 57334 321600
rect 57390 321558 60076 321600
rect 57390 321544 59554 321558
rect 57329 321542 59554 321544
rect 57329 321539 57395 321542
rect 406653 320786 406719 320789
rect 404678 320784 406719 320786
rect 404678 320762 406658 320784
rect 404064 320728 406658 320762
rect 406714 320728 406719 320784
rect 404064 320726 406719 320728
rect 404064 320702 404738 320726
rect 406653 320723 406719 320726
rect -960 319290 480 319380
rect 3141 319290 3207 319293
rect -960 319288 3207 319290
rect -960 319232 3146 319288
rect 3202 319232 3207 319288
rect -960 319230 3207 319232
rect -960 319140 480 319230
rect 3141 319227 3207 319230
rect 57605 316162 57671 316165
rect 57605 316160 59554 316162
rect 57605 316104 57610 316160
rect 57666 316104 59554 316160
rect 57605 316102 59554 316104
rect 57605 316099 57671 316102
rect 59494 316072 59554 316102
rect 59494 316012 60076 316072
rect 404064 315074 404738 315109
rect 406745 315074 406811 315077
rect 404064 315072 406811 315074
rect 404064 315049 406750 315072
rect 404678 315016 406750 315049
rect 406806 315016 406811 315072
rect 404678 315014 406811 315016
rect 406745 315011 406811 315014
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 59494 310465 60076 310525
rect 57605 310450 57671 310453
rect 59494 310450 59554 310465
rect 57605 310448 59554 310450
rect 57605 310392 57610 310448
rect 57666 310392 59554 310448
rect 57605 310390 59554 310392
rect 57605 310387 57671 310390
rect 406837 309498 406903 309501
rect 404678 309496 406903 309498
rect 404678 309456 406842 309496
rect 404064 309440 406842 309456
rect 406898 309440 406903 309496
rect 404064 309438 406903 309440
rect 404064 309396 404738 309438
rect 406837 309435 406903 309438
rect -960 306234 480 306324
rect 3049 306234 3115 306237
rect -960 306232 3115 306234
rect -960 306176 3054 306232
rect 3110 306176 3115 306232
rect -960 306174 3115 306176
rect -960 306084 480 306174
rect 3049 306171 3115 306174
rect 57421 305010 57487 305013
rect 57421 305008 59554 305010
rect 57421 304952 57426 305008
rect 57482 304979 59554 305008
rect 57482 304952 60076 304979
rect 57421 304950 60076 304952
rect 57421 304947 57487 304950
rect 59494 304919 60076 304950
rect 404064 303786 404738 303803
rect 406837 303786 406903 303789
rect 404064 303784 406903 303786
rect 404064 303743 406842 303784
rect 404678 303728 406842 303743
rect 406898 303728 406903 303784
rect 404678 303726 406903 303728
rect 406837 303723 406903 303726
rect 57605 299434 57671 299437
rect 57605 299432 59554 299434
rect 57605 299376 57610 299432
rect 57666 299376 60076 299432
rect 57605 299374 60076 299376
rect 57605 299371 57671 299374
rect 59494 299372 60076 299374
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 405825 298210 405891 298213
rect 404678 298208 405891 298210
rect 404678 298152 405830 298208
rect 405886 298152 405891 298208
rect 404678 298150 405891 298152
rect 404064 298090 404738 298150
rect 405825 298147 405891 298150
rect 57605 293858 57671 293861
rect 59494 293858 60076 293886
rect 57605 293856 60076 293858
rect 57605 293800 57610 293856
rect 57666 293826 60076 293856
rect 57666 293800 59554 293826
rect 57605 293798 59554 293800
rect 57605 293795 57671 293798
rect -960 293178 480 293268
rect 2957 293178 3023 293181
rect -960 293176 3023 293178
rect -960 293120 2962 293176
rect 3018 293120 3023 293176
rect -960 293118 3023 293120
rect -960 293028 480 293118
rect 2957 293115 3023 293118
rect 406837 292498 406903 292501
rect 404678 292497 406903 292498
rect 404064 292496 406903 292497
rect 404064 292440 406842 292496
rect 406898 292440 406903 292496
rect 404064 292438 406903 292440
rect 404064 292437 404738 292438
rect 406837 292435 406903 292438
rect 57605 288418 57671 288421
rect 57605 288416 59554 288418
rect 57605 288360 57610 288416
rect 57666 288360 59554 288416
rect 57605 288358 59554 288360
rect 57605 288355 57671 288358
rect 59494 288340 59554 288358
rect 59494 288280 60076 288340
rect 404064 286786 404738 286844
rect 406837 286786 406903 286789
rect 404064 286784 406903 286786
rect 404678 286728 406842 286784
rect 406898 286728 406903 286784
rect 404678 286726 406903 286728
rect 406837 286723 406903 286726
rect 580349 285426 580415 285429
rect 583520 285426 584960 285516
rect 580349 285424 584960 285426
rect 580349 285368 580354 285424
rect 580410 285368 584960 285424
rect 580349 285366 584960 285368
rect 580349 285363 580415 285366
rect 583520 285276 584960 285366
rect 57605 282842 57671 282845
rect 57605 282840 59554 282842
rect 57605 282784 57610 282840
rect 57666 282793 59554 282840
rect 57666 282784 60076 282793
rect 57605 282782 60076 282784
rect 57605 282779 57671 282782
rect 59494 282733 60076 282782
rect 406837 281210 406903 281213
rect 404678 281208 406903 281210
rect 404678 281191 406842 281208
rect 404064 281152 406842 281191
rect 406898 281152 406903 281208
rect 404064 281150 406903 281152
rect 404064 281131 404738 281150
rect 406837 281147 406903 281150
rect -960 280122 480 280212
rect 3693 280122 3759 280125
rect -960 280120 3759 280122
rect -960 280064 3698 280120
rect 3754 280064 3759 280120
rect -960 280062 3759 280064
rect -960 279972 480 280062
rect 3693 280059 3759 280062
rect 57605 277266 57671 277269
rect 57605 277264 59554 277266
rect 57605 277208 57610 277264
rect 57666 277247 59554 277264
rect 57666 277208 60076 277247
rect 57605 277206 60076 277208
rect 57605 277203 57671 277206
rect 59494 277187 60076 277206
rect 404064 275498 404738 275538
rect 406929 275498 406995 275501
rect 404064 275496 406995 275498
rect 404064 275478 406934 275496
rect 404678 275440 406934 275478
rect 406990 275440 406995 275496
rect 404678 275438 406995 275440
rect 406929 275435 406995 275438
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 57513 271690 57579 271693
rect 59494 271690 60076 271700
rect 57513 271688 60076 271690
rect 57513 271632 57518 271688
rect 57574 271640 60076 271688
rect 57574 271632 59554 271640
rect 57513 271630 59554 271632
rect 57513 271627 57579 271630
rect 407021 269922 407087 269925
rect 404678 269920 407087 269922
rect 404678 269885 407026 269920
rect 404064 269864 407026 269885
rect 407082 269864 407087 269920
rect 404064 269862 407087 269864
rect 404064 269825 404738 269862
rect 407021 269859 407087 269862
rect -960 267202 480 267292
rect 3785 267202 3851 267205
rect -960 267200 3851 267202
rect -960 267144 3790 267200
rect 3846 267144 3851 267200
rect -960 267142 3851 267144
rect -960 267052 480 267142
rect 3785 267139 3851 267142
rect 57329 266114 57395 266117
rect 59494 266114 60076 266154
rect 57329 266112 60076 266114
rect 57329 266056 57334 266112
rect 57390 266094 60076 266112
rect 57390 266056 59554 266094
rect 57329 266054 59554 266056
rect 57329 266051 57395 266054
rect 404064 264210 404738 264232
rect 407021 264210 407087 264213
rect 404064 264208 407087 264210
rect 404064 264172 407026 264208
rect 404678 264152 407026 264172
rect 407082 264152 407087 264208
rect 404678 264150 407087 264152
rect 407021 264147 407087 264150
rect 57421 260674 57487 260677
rect 57421 260672 59554 260674
rect 57421 260616 57426 260672
rect 57482 260616 59554 260672
rect 57421 260614 59554 260616
rect 57421 260611 57487 260614
rect 59494 260608 59554 260614
rect 59494 260548 60076 260608
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 404064 258519 404738 258579
rect 404678 257954 404738 258519
rect 406929 258090 406995 258093
rect 406886 258088 406995 258090
rect 406886 258032 406934 258088
rect 406990 258032 406995 258088
rect 406886 258027 406995 258032
rect 406886 257954 406946 258027
rect 404678 257894 406946 257954
rect 57605 255098 57671 255101
rect 57605 255096 59554 255098
rect 57605 255040 57610 255096
rect 57666 255061 59554 255096
rect 57666 255040 60076 255061
rect 57605 255038 60076 255040
rect 57605 255035 57671 255038
rect 59494 255001 60076 255038
rect -960 254146 480 254236
rect 2865 254146 2931 254149
rect -960 254144 2931 254146
rect -960 254088 2870 254144
rect 2926 254088 2931 254144
rect -960 254086 2931 254088
rect -960 253996 480 254086
rect 2865 254083 2931 254086
rect 404064 252922 404738 252926
rect 407021 252922 407087 252925
rect 404064 252920 407087 252922
rect 404064 252866 407026 252920
rect 404678 252864 407026 252866
rect 407082 252864 407087 252920
rect 404678 252862 407087 252864
rect 407021 252859 407087 252862
rect 57237 249522 57303 249525
rect 57237 249520 59554 249522
rect 57237 249464 57242 249520
rect 57298 249515 59554 249520
rect 57298 249464 60076 249515
rect 57237 249462 60076 249464
rect 57237 249459 57303 249462
rect 59494 249455 60076 249462
rect 404064 247213 404738 247273
rect 404678 247210 404738 247213
rect 406285 247210 406351 247213
rect 404678 247208 406351 247210
rect 404678 247152 406290 247208
rect 406346 247152 406351 247208
rect 404678 247150 406351 247152
rect 406285 247147 406351 247150
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 57421 243946 57487 243949
rect 59494 243946 60076 243968
rect 57421 243944 60076 243946
rect 57421 243888 57426 243944
rect 57482 243908 60076 243944
rect 57482 243888 59554 243908
rect 57421 243886 59554 243888
rect 57421 243883 57487 243886
rect 406193 241634 406259 241637
rect 404678 241632 406259 241634
rect 404678 241620 406198 241632
rect 404064 241576 406198 241620
rect 406254 241576 406259 241632
rect 404064 241574 406259 241576
rect 404064 241560 404738 241574
rect 406193 241571 406259 241574
rect -960 241090 480 241180
rect 3877 241090 3943 241093
rect -960 241088 3943 241090
rect -960 241032 3882 241088
rect 3938 241032 3943 241088
rect -960 241030 3943 241032
rect -960 240940 480 241030
rect 3877 241027 3943 241030
rect 57605 238506 57671 238509
rect 57605 238504 59554 238506
rect 57605 238448 57610 238504
rect 57666 238448 59554 238504
rect 57605 238446 59554 238448
rect 57605 238443 57671 238446
rect 59494 238422 59554 238446
rect 59494 238362 60076 238422
rect 404064 235922 404738 235967
rect 407021 235922 407087 235925
rect 404064 235920 407087 235922
rect 404064 235907 407026 235920
rect 404678 235864 407026 235907
rect 407082 235864 407087 235920
rect 404678 235862 407087 235864
rect 407021 235859 407087 235862
rect 57605 232930 57671 232933
rect 57605 232928 59554 232930
rect 57605 232872 57610 232928
rect 57666 232876 59554 232928
rect 57666 232872 60076 232876
rect 57605 232870 60076 232872
rect 57605 232867 57671 232870
rect 59494 232816 60076 232870
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect 406101 230346 406167 230349
rect 404678 230344 406167 230346
rect 404678 230314 406106 230344
rect 404064 230288 406106 230314
rect 406162 230288 406167 230344
rect 404064 230286 406167 230288
rect 404064 230254 404738 230286
rect 406101 230283 406167 230286
rect -960 228034 480 228124
rect 3969 228034 4035 228037
rect -960 228032 4035 228034
rect -960 227976 3974 228032
rect 4030 227976 4035 228032
rect -960 227974 4035 227976
rect -960 227884 480 227974
rect 3969 227971 4035 227974
rect 57605 227354 57671 227357
rect 57605 227352 59554 227354
rect 57605 227296 57610 227352
rect 57666 227329 59554 227352
rect 57666 227296 60076 227329
rect 57605 227294 60076 227296
rect 57605 227291 57671 227294
rect 59494 227269 60076 227294
rect 404064 224634 404738 224661
rect 406285 224634 406351 224637
rect 404064 224632 406351 224634
rect 404064 224601 406290 224632
rect 404678 224576 406290 224601
rect 406346 224576 406351 224632
rect 404678 224574 406351 224576
rect 406285 224571 406351 224574
rect 57605 221778 57671 221781
rect 59494 221778 60076 221783
rect 57605 221776 60076 221778
rect 57605 221720 57610 221776
rect 57666 221723 60076 221776
rect 57666 221720 59554 221723
rect 57605 221718 59554 221720
rect 57605 221715 57671 221718
rect 406377 219058 406443 219061
rect 404678 219056 406443 219058
rect 404678 219008 406382 219056
rect 404064 219000 406382 219008
rect 406438 219000 406443 219056
rect 404064 218998 406443 219000
rect 404064 218948 404738 218998
rect 406377 218995 406443 218998
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 57053 216202 57119 216205
rect 59494 216202 60076 216236
rect 57053 216200 60076 216202
rect 57053 216144 57058 216200
rect 57114 216176 60076 216200
rect 57114 216144 59554 216176
rect 57053 216142 59554 216144
rect 57053 216139 57119 216142
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 404064 213346 404738 213355
rect 406377 213346 406443 213349
rect 404064 213344 406443 213346
rect 404064 213295 406382 213344
rect 404678 213288 406382 213295
rect 406438 213288 406443 213344
rect 404678 213286 406443 213288
rect 406377 213283 406443 213286
rect 56777 210762 56843 210765
rect 56777 210760 59554 210762
rect 56777 210704 56782 210760
rect 56838 210704 59554 210760
rect 56777 210702 59554 210704
rect 56777 210699 56843 210702
rect 59494 210690 59554 210702
rect 59494 210630 60076 210690
rect 406469 207770 406535 207773
rect 404310 207768 406535 207770
rect 404310 207712 406474 207768
rect 406530 207712 406535 207768
rect 404310 207710 406535 207712
rect 404310 207702 404370 207710
rect 406469 207707 406535 207710
rect 404064 207642 404370 207702
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 57605 205186 57671 205189
rect 57605 205184 59554 205186
rect 57605 205128 57610 205184
rect 57666 205144 59554 205184
rect 57666 205128 60076 205144
rect 57605 205126 60076 205128
rect 57605 205123 57671 205126
rect 59494 205084 60076 205126
rect 406561 202058 406627 202061
rect 404678 202056 406627 202058
rect 404678 202049 406566 202056
rect -960 201922 480 202012
rect 404064 202000 406566 202049
rect 406622 202000 406627 202056
rect 404064 201998 406627 202000
rect 404064 201989 404738 201998
rect 406561 201995 406627 201998
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 57605 199610 57671 199613
rect 57605 199608 59554 199610
rect 57605 199552 57610 199608
rect 57666 199597 59554 199608
rect 57666 199552 60076 199597
rect 57605 199550 60076 199552
rect 57605 199547 57671 199550
rect 59494 199537 60076 199550
rect 404064 196346 404738 196396
rect 406653 196346 406719 196349
rect 404064 196344 406719 196346
rect 404064 196336 406658 196344
rect 404678 196288 406658 196336
rect 406714 196288 406719 196344
rect 404678 196286 406719 196288
rect 406653 196283 406719 196286
rect 57605 194034 57671 194037
rect 59494 194034 60076 194051
rect 57605 194032 60076 194034
rect 57605 193976 57610 194032
rect 57666 193991 60076 194032
rect 57666 193976 59554 193991
rect 57605 193974 59554 193976
rect 57605 193971 57671 193974
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 406745 190770 406811 190773
rect 404678 190768 406811 190770
rect 404678 190743 406750 190768
rect 404064 190712 406750 190743
rect 406806 190712 406811 190768
rect 404064 190710 406811 190712
rect 404064 190683 404738 190710
rect 406745 190707 406811 190710
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 57605 188594 57671 188597
rect 57605 188592 59554 188594
rect 57605 188536 57610 188592
rect 57666 188536 59554 188592
rect 57605 188534 59554 188536
rect 57605 188531 57671 188534
rect 59494 188504 59554 188534
rect 59494 188444 60076 188504
rect 404064 185058 404738 185090
rect 406653 185058 406719 185061
rect 404064 185056 406719 185058
rect 404064 185030 406658 185056
rect 404678 185000 406658 185030
rect 406714 185000 406719 185056
rect 404678 184998 406719 185000
rect 406653 184995 406719 184998
rect 57605 183018 57671 183021
rect 57605 183016 59554 183018
rect 57605 182960 57610 183016
rect 57666 182960 59554 183016
rect 57605 182958 59554 182960
rect 57605 182955 57671 182958
rect 59494 182898 60076 182958
rect 406837 179482 406903 179485
rect 404678 179480 406903 179482
rect 404678 179437 406842 179480
rect 404064 179424 406842 179437
rect 406898 179424 406903 179480
rect 404064 179422 406903 179424
rect 404064 179377 404738 179422
rect 406837 179419 406903 179422
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 56685 177442 56751 177445
rect 56685 177440 59554 177442
rect 56685 177384 56690 177440
rect 56746 177412 59554 177440
rect 56746 177384 60076 177412
rect 56685 177382 60076 177384
rect 56685 177379 56751 177382
rect 59494 177352 60076 177382
rect -960 175946 480 176036
rect 3693 175946 3759 175949
rect -960 175944 3759 175946
rect -960 175888 3698 175944
rect 3754 175888 3759 175944
rect -960 175886 3759 175888
rect -960 175796 480 175886
rect 3693 175883 3759 175886
rect 404064 173770 404738 173784
rect 406929 173770 406995 173773
rect 404064 173768 406995 173770
rect 404064 173724 406934 173768
rect 404678 173712 406934 173724
rect 406990 173712 406995 173768
rect 404678 173710 406995 173712
rect 406929 173707 406995 173710
rect 57605 171866 57671 171869
rect 57605 171865 59554 171866
rect 57605 171864 60076 171865
rect 57605 171808 57610 171864
rect 57666 171808 60076 171864
rect 57605 171806 60076 171808
rect 57605 171803 57671 171806
rect 59494 171805 60076 171806
rect 407021 168194 407087 168197
rect 404678 168192 407087 168194
rect 404678 168136 407026 168192
rect 407082 168136 407087 168192
rect 404678 168134 407087 168136
rect 404678 168131 404738 168134
rect 407021 168131 407087 168134
rect 404064 168071 404738 168131
rect 57605 166290 57671 166293
rect 59494 166290 60076 166319
rect 57605 166288 60076 166290
rect 57605 166232 57610 166288
rect 57666 166259 60076 166288
rect 57666 166232 59554 166259
rect 57605 166230 59554 166232
rect 57605 166227 57671 166230
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3785 162890 3851 162893
rect -960 162888 3851 162890
rect -960 162832 3790 162888
rect 3846 162832 3851 162888
rect -960 162830 3851 162832
rect -960 162740 480 162830
rect 3785 162827 3851 162830
rect 406285 162482 406351 162485
rect 404678 162480 406351 162482
rect 404678 162478 406290 162480
rect 404064 162424 406290 162478
rect 406346 162424 406351 162480
rect 404064 162422 406351 162424
rect 404064 162418 404738 162422
rect 406285 162419 406351 162422
rect 57605 160850 57671 160853
rect 57605 160848 59554 160850
rect 57605 160792 57610 160848
rect 57666 160792 59554 160848
rect 57605 160790 59554 160792
rect 57605 160787 57671 160790
rect 59494 160772 59554 160790
rect 59494 160712 60076 160772
rect 404064 156770 404738 156825
rect 406377 156770 406443 156773
rect 404064 156768 406443 156770
rect 404064 156765 406382 156768
rect 404678 156712 406382 156765
rect 406438 156712 406443 156768
rect 404678 156710 406443 156712
rect 406377 156707 406443 156710
rect 57605 155274 57671 155277
rect 57605 155272 59554 155274
rect 57605 155216 57610 155272
rect 57666 155226 59554 155272
rect 57666 155216 60076 155226
rect 57605 155214 60076 155216
rect 57605 155211 57671 155214
rect 59494 155166 60076 155214
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect 406469 151194 406535 151197
rect 404678 151192 406535 151194
rect 404678 151172 406474 151192
rect 404064 151136 406474 151172
rect 406530 151136 406535 151192
rect 404064 151134 406535 151136
rect 404064 151112 404738 151134
rect 406469 151131 406535 151134
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 56869 149698 56935 149701
rect 56869 149696 59554 149698
rect 56869 149640 56874 149696
rect 56930 149680 59554 149696
rect 56930 149640 60076 149680
rect 56869 149638 60076 149640
rect 56869 149635 56935 149638
rect 59494 149620 60076 149638
rect 404064 145482 404738 145519
rect 406561 145482 406627 145485
rect 404064 145480 406627 145482
rect 404064 145459 406566 145480
rect 404678 145424 406566 145459
rect 406622 145424 406627 145480
rect 404678 145422 406627 145424
rect 406561 145419 406627 145422
rect 57513 144122 57579 144125
rect 59494 144122 60076 144133
rect 57513 144120 60076 144122
rect 57513 144064 57518 144120
rect 57574 144073 60076 144120
rect 57574 144064 59554 144073
rect 57513 144062 59554 144064
rect 57513 144059 57579 144062
rect 406653 139906 406719 139909
rect 404678 139904 406719 139906
rect 404678 139866 406658 139904
rect 404064 139848 406658 139866
rect 406714 139848 406719 139904
rect 404064 139846 406719 139848
rect 404064 139806 404738 139846
rect 406653 139843 406719 139846
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 57513 138546 57579 138549
rect 59494 138546 60076 138587
rect 57513 138544 60076 138546
rect 57513 138488 57518 138544
rect 57574 138527 60076 138544
rect 57574 138488 59554 138527
rect 57513 138486 59554 138488
rect 57513 138483 57579 138486
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 404064 134194 404738 134213
rect 406377 134194 406443 134197
rect 404064 134192 406443 134194
rect 404064 134153 406382 134192
rect 404678 134136 406382 134153
rect 406438 134136 406443 134192
rect 404678 134134 406443 134136
rect 406377 134131 406443 134134
rect 57513 133106 57579 133109
rect 57513 133104 59554 133106
rect 57513 133048 57518 133104
rect 57574 133048 59554 133104
rect 57513 133046 59554 133048
rect 57513 133043 57579 133046
rect 59494 133040 59554 133046
rect 59494 132980 60076 133040
rect 406469 128618 406535 128621
rect 404678 128616 406535 128618
rect 404678 128560 406474 128616
rect 406530 128560 406535 128616
rect 404064 128558 406535 128560
rect 404064 128500 404738 128558
rect 406469 128555 406535 128558
rect 56961 127530 57027 127533
rect 56961 127528 59554 127530
rect 56961 127472 56966 127528
rect 57022 127494 59554 127528
rect 57022 127472 60076 127494
rect 56961 127470 60076 127472
rect 56961 127467 57027 127470
rect 59494 127434 60076 127470
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 3601 123722 3667 123725
rect -960 123720 3667 123722
rect -960 123664 3606 123720
rect 3662 123664 3667 123720
rect -960 123662 3667 123664
rect -960 123572 480 123662
rect 3601 123659 3667 123662
rect 404064 122906 404738 122907
rect 407021 122906 407087 122909
rect 404064 122904 407087 122906
rect 404064 122848 407026 122904
rect 407082 122848 407087 122904
rect 404064 122847 407087 122848
rect 404678 122846 407087 122847
rect 407021 122843 407087 122846
rect 57053 121954 57119 121957
rect 57053 121952 59554 121954
rect 57053 121896 57058 121952
rect 57114 121948 59554 121952
rect 57114 121896 60076 121948
rect 57053 121894 60076 121896
rect 57053 121891 57119 121894
rect 59494 121888 60076 121894
rect 404064 117194 404738 117254
rect 406377 117194 406443 117197
rect 404678 117192 406443 117194
rect 404678 117136 406382 117192
rect 406438 117136 406443 117192
rect 404678 117134 406443 117136
rect 406377 117131 406443 117134
rect 57605 116378 57671 116381
rect 59494 116378 60076 116401
rect 57605 116376 60076 116378
rect 57605 116320 57610 116376
rect 57666 116341 60076 116376
rect 57666 116320 59554 116341
rect 57605 116318 59554 116320
rect 57605 116315 57671 116318
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 406469 111618 406535 111621
rect 404678 111616 406535 111618
rect 404678 111601 406474 111616
rect 404064 111560 406474 111601
rect 406530 111560 406535 111616
rect 404064 111558 406535 111560
rect 404064 111541 404738 111558
rect 406469 111555 406535 111558
rect 57605 110802 57671 110805
rect 59494 110802 60076 110855
rect 57605 110800 60076 110802
rect -960 110666 480 110756
rect 57605 110744 57610 110800
rect 57666 110795 60076 110800
rect 57666 110744 59554 110795
rect 57605 110742 59554 110744
rect 57605 110739 57671 110742
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 404064 105906 404738 105948
rect 406377 105906 406443 105909
rect 404064 105904 406443 105906
rect 404064 105888 406382 105904
rect 404678 105848 406382 105888
rect 406438 105848 406443 105904
rect 404678 105846 406443 105848
rect 406377 105843 406443 105846
rect 59494 105248 60076 105308
rect 57421 105226 57487 105229
rect 59494 105226 59554 105248
rect 57421 105224 59554 105226
rect 57421 105168 57426 105224
rect 57482 105168 59554 105224
rect 57421 105166 59554 105168
rect 57421 105163 57487 105166
rect 406837 100330 406903 100333
rect 404678 100328 406903 100330
rect 404678 100295 406842 100328
rect 404064 100272 406842 100295
rect 406898 100272 406903 100328
rect 404064 100270 406903 100272
rect 404064 100235 404738 100270
rect 406837 100267 406903 100270
rect 57421 99786 57487 99789
rect 57421 99784 59554 99786
rect 57421 99728 57426 99784
rect 57482 99762 59554 99784
rect 57482 99728 60076 99762
rect 57421 99726 60076 99728
rect 57421 99723 57487 99726
rect 59494 99702 60076 99726
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 404064 94618 404738 94642
rect 406745 94618 406811 94621
rect 404064 94616 406811 94618
rect 404064 94582 406750 94616
rect 404678 94560 406750 94582
rect 406806 94560 406811 94616
rect 404678 94558 406811 94560
rect 406745 94555 406811 94558
rect 57605 94210 57671 94213
rect 59494 94210 60076 94216
rect 57605 94208 60076 94210
rect 57605 94152 57610 94208
rect 57666 94156 60076 94208
rect 57666 94152 59554 94156
rect 57605 94150 59554 94152
rect 57605 94147 57671 94150
rect 404064 88929 404738 88989
rect 404678 88906 404738 88929
rect 406653 88906 406719 88909
rect 404678 88904 406719 88906
rect 404678 88848 406658 88904
rect 406714 88848 406719 88904
rect 404678 88846 406719 88848
rect 406653 88843 406719 88846
rect 57513 88634 57579 88637
rect 59494 88634 60076 88669
rect 57513 88632 60076 88634
rect 57513 88576 57518 88632
rect 57574 88609 60076 88632
rect 57574 88576 59554 88609
rect 57513 88574 59554 88576
rect 57513 88571 57579 88574
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 404064 83330 404738 83336
rect 406561 83330 406627 83333
rect 404064 83328 406627 83330
rect 404064 83276 406566 83328
rect 404678 83272 406566 83276
rect 406622 83272 406627 83328
rect 404678 83270 406627 83272
rect 406561 83267 406627 83270
rect 59494 83063 60076 83123
rect 57421 83058 57487 83061
rect 59494 83058 59554 83063
rect 57421 83056 59554 83058
rect 57421 83000 57426 83056
rect 57482 83000 59554 83056
rect 57421 82998 59554 83000
rect 57421 82995 57487 82998
rect 404064 77623 404738 77683
rect 57513 77618 57579 77621
rect 404678 77618 404738 77623
rect 406469 77618 406535 77621
rect 57513 77616 59554 77618
rect 57513 77560 57518 77616
rect 57574 77576 59554 77616
rect 404678 77616 406535 77618
rect 57574 77560 60076 77576
rect 57513 77558 60076 77560
rect 404678 77560 406474 77616
rect 406530 77560 406535 77616
rect 404678 77558 406535 77560
rect 57513 77555 57579 77558
rect 59494 77516 60076 77558
rect 406469 77555 406535 77558
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 59494 72878 60076 72938
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 57421 72858 57487 72861
rect 59494 72858 59554 72878
rect 406377 72858 406443 72861
rect 57421 72856 59554 72858
rect 57421 72800 57426 72856
rect 57482 72800 59554 72856
rect 404678 72856 406443 72858
rect 404678 72816 406382 72856
rect 57421 72798 59554 72800
rect 404064 72800 406382 72816
rect 406438 72800 406443 72856
rect 583520 72844 584960 72934
rect 404064 72798 406443 72800
rect 57421 72795 57487 72798
rect 404064 72756 404738 72798
rect 406377 72795 406443 72798
rect -960 71634 480 71724
rect 3877 71634 3943 71637
rect -960 71632 3943 71634
rect -960 71576 3882 71632
rect 3938 71576 3943 71632
rect -960 71574 3943 71576
rect -960 71484 480 71574
rect 3877 71571 3943 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3785 58578 3851 58581
rect -960 58576 3851 58578
rect -960 58520 3790 58576
rect 3846 58520 3851 58576
rect -960 58518 3851 58520
rect -960 58428 480 58518
rect 3785 58515 3851 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3693 45522 3759 45525
rect -960 45520 3759 45522
rect -960 45464 3698 45520
rect 3754 45464 3759 45520
rect -960 45462 3759 45464
rect -960 45372 480 45462
rect 3693 45459 3759 45462
rect 579889 33146 579955 33149
rect 583520 33146 584960 33236
rect 579889 33144 584960 33146
rect 579889 33088 579894 33144
rect 579950 33088 584960 33144
rect 579889 33086 584960 33088
rect 579889 33083 579955 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3601 32466 3667 32469
rect -960 32464 3667 32466
rect -960 32408 3606 32464
rect 3662 32408 3667 32464
rect -960 32406 3667 32408
rect -960 32316 480 32406
rect 3601 32403 3667 32406
rect 579889 19818 579955 19821
rect 583520 19818 584960 19908
rect 579889 19816 584960 19818
rect 579889 19760 579894 19816
rect 579950 19760 584960 19816
rect 579889 19758 584960 19760
rect 579889 19755 579955 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 25313 3770 25379 3773
rect 131205 3770 131271 3773
rect 25313 3768 131271 3770
rect 25313 3712 25318 3768
rect 25374 3712 131210 3768
rect 131266 3712 131271 3768
rect 25313 3710 131271 3712
rect 25313 3707 25379 3710
rect 131205 3707 131271 3710
rect 245193 3770 245259 3773
rect 335537 3770 335603 3773
rect 245193 3768 335603 3770
rect 245193 3712 245198 3768
rect 245254 3712 335542 3768
rect 335598 3712 335603 3768
rect 245193 3710 335603 3712
rect 245193 3707 245259 3710
rect 335537 3707 335603 3710
rect 404261 3770 404327 3773
rect 582189 3770 582255 3773
rect 404261 3768 582255 3770
rect 404261 3712 404266 3768
rect 404322 3712 582194 3768
rect 582250 3712 582255 3768
rect 404261 3710 582255 3712
rect 404261 3707 404327 3710
rect 582189 3707 582255 3710
rect 20621 3634 20687 3637
rect 131113 3634 131179 3637
rect 20621 3632 131179 3634
rect 20621 3576 20626 3632
rect 20682 3576 131118 3632
rect 131174 3576 131179 3632
rect 20621 3574 131179 3576
rect 20621 3571 20687 3574
rect 131113 3571 131179 3574
rect 241697 3634 241763 3637
rect 333973 3634 334039 3637
rect 241697 3632 334039 3634
rect 241697 3576 241702 3632
rect 241758 3576 333978 3632
rect 334034 3576 334039 3632
rect 241697 3574 334039 3576
rect 241697 3571 241763 3574
rect 333973 3571 334039 3574
rect 401409 3634 401475 3637
rect 578601 3634 578667 3637
rect 401409 3632 578667 3634
rect 401409 3576 401414 3632
rect 401470 3576 578606 3632
rect 578662 3576 578667 3632
rect 401409 3574 578667 3576
rect 401409 3571 401475 3574
rect 578601 3571 578667 3574
rect 11145 3498 11211 3501
rect 129825 3498 129891 3501
rect 11145 3496 129891 3498
rect 11145 3440 11150 3496
rect 11206 3440 129830 3496
rect 129886 3440 129891 3496
rect 11145 3438 129891 3440
rect 11145 3435 11211 3438
rect 129825 3435 129891 3438
rect 142429 3498 142495 3501
rect 314745 3498 314811 3501
rect 142429 3496 314811 3498
rect 142429 3440 142434 3496
rect 142490 3440 314750 3496
rect 314806 3440 314811 3496
rect 142429 3438 314811 3440
rect 142429 3435 142495 3438
rect 314745 3435 314811 3438
rect 402789 3498 402855 3501
rect 580993 3498 581059 3501
rect 402789 3496 581059 3498
rect 402789 3440 402794 3496
rect 402850 3440 580998 3496
rect 581054 3440 581059 3496
rect 402789 3438 581059 3440
rect 402789 3435 402855 3438
rect 580993 3435 581059 3438
rect 5257 3362 5323 3365
rect 132585 3362 132651 3365
rect 5257 3360 132651 3362
rect 5257 3304 5262 3360
rect 5318 3304 132590 3360
rect 132646 3304 132651 3360
rect 5257 3302 132651 3304
rect 5257 3299 5323 3302
rect 132585 3299 132651 3302
rect 138841 3362 138907 3365
rect 314837 3362 314903 3365
rect 138841 3360 314903 3362
rect 138841 3304 138846 3360
rect 138902 3304 314842 3360
rect 314898 3304 314903 3360
rect 138841 3302 314903 3304
rect 138841 3299 138907 3302
rect 314837 3299 314903 3302
rect 402881 3362 402947 3365
rect 583385 3362 583451 3365
rect 402881 3360 583451 3362
rect 402881 3304 402886 3360
rect 402942 3304 583390 3360
rect 583446 3304 583451 3360
rect 402881 3302 583451 3304
rect 402881 3299 402947 3302
rect 583385 3299 583451 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 367964 60134 384618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 367964 63854 388338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 367964 67574 392058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 367964 74414 398898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367964 78134 402618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 367964 81854 370338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 367964 85574 374058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 367964 92414 380898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 367964 96134 384618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 367964 99854 388338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 367964 103574 392058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 367964 110414 398898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367964 114134 402618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 367964 117854 370338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 367964 121574 374058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 367964 128414 380898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 367964 132134 384618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 367964 135854 388338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 367964 139574 392058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 367964 146414 398898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367964 150134 402618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 367964 153854 370338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 367964 157574 374058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 367964 164414 380898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 367964 168134 384618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 367964 171854 388338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 367964 175574 392058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 367964 182414 398898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367964 186134 402618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 367964 189854 370338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 367964 193574 374058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 367964 200414 380898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 367964 204134 384618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 367964 207854 388338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 367964 211574 392058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 367964 218414 398898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367964 222134 402618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 367964 225854 370338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 367964 229574 374058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 367964 236414 380898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 367964 240134 384618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 367964 243854 388338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 367964 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 367964 254414 398898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367964 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 367964 261854 370338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 367964 265574 374058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 367964 272414 380898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 367964 276134 384618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 367964 279854 388338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 367964 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 367964 290414 398898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367964 294134 402618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 367964 297854 370338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 367964 301574 374058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 367964 308414 380898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 367964 312134 384618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 367964 315854 388338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 367964 319574 392058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 367964 326414 398898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367964 330134 402618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 367964 333854 370338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 367964 337574 374058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 367964 344414 380898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 367964 348134 384618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 367964 351854 388338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 367964 355574 392058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 367964 362414 398898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367964 366134 402618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 367964 369854 370338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 367964 373574 374058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 367964 380414 380898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 367964 384134 384618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 367964 387854 388338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 367964 391574 392058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 367964 398414 398898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367964 402134 402618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 367964 405854 370338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 60412 363454 60812 363486
rect 60412 363218 60494 363454
rect 60730 363218 60812 363454
rect 60412 363134 60812 363218
rect 60412 362898 60494 363134
rect 60730 362898 60812 363134
rect 60412 362866 60812 362898
rect 403268 363454 403668 363486
rect 403268 363218 403350 363454
rect 403586 363218 403668 363454
rect 403268 363134 403668 363218
rect 403268 362898 403350 363134
rect 403586 362898 403668 363134
rect 403268 362866 403668 362898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 61212 345454 61612 345486
rect 61212 345218 61294 345454
rect 61530 345218 61612 345454
rect 61212 345134 61612 345218
rect 61212 344898 61294 345134
rect 61530 344898 61612 345134
rect 61212 344866 61612 344898
rect 402468 345454 402868 345486
rect 402468 345218 402550 345454
rect 402786 345218 402868 345454
rect 402468 345134 402868 345218
rect 402468 344898 402550 345134
rect 402786 344898 402868 345134
rect 402468 344866 402868 344898
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 60412 327454 60812 327486
rect 60412 327218 60494 327454
rect 60730 327218 60812 327454
rect 60412 327134 60812 327218
rect 60412 326898 60494 327134
rect 60730 326898 60812 327134
rect 60412 326866 60812 326898
rect 403268 327454 403668 327486
rect 403268 327218 403350 327454
rect 403586 327218 403668 327454
rect 403268 327134 403668 327218
rect 403268 326898 403350 327134
rect 403586 326898 403668 327134
rect 403268 326866 403668 326898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 61212 309454 61612 309486
rect 61212 309218 61294 309454
rect 61530 309218 61612 309454
rect 61212 309134 61612 309218
rect 61212 308898 61294 309134
rect 61530 308898 61612 309134
rect 61212 308866 61612 308898
rect 402468 309454 402868 309486
rect 402468 309218 402550 309454
rect 402786 309218 402868 309454
rect 402468 309134 402868 309218
rect 402468 308898 402550 309134
rect 402786 308898 402868 309134
rect 402468 308866 402868 308898
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 60412 291454 60812 291486
rect 60412 291218 60494 291454
rect 60730 291218 60812 291454
rect 60412 291134 60812 291218
rect 60412 290898 60494 291134
rect 60730 290898 60812 291134
rect 60412 290866 60812 290898
rect 403268 291454 403668 291486
rect 403268 291218 403350 291454
rect 403586 291218 403668 291454
rect 403268 291134 403668 291218
rect 403268 290898 403350 291134
rect 403586 290898 403668 291134
rect 403268 290866 403668 290898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 61212 273454 61612 273486
rect 61212 273218 61294 273454
rect 61530 273218 61612 273454
rect 61212 273134 61612 273218
rect 61212 272898 61294 273134
rect 61530 272898 61612 273134
rect 61212 272866 61612 272898
rect 77013 273454 77361 273486
rect 77013 273218 77069 273454
rect 77305 273218 77361 273454
rect 77013 273134 77361 273218
rect 77013 272898 77069 273134
rect 77305 272898 77361 273134
rect 77013 272866 77361 272898
rect 172077 273454 172425 273486
rect 172077 273218 172133 273454
rect 172369 273218 172425 273454
rect 172077 273134 172425 273218
rect 172077 272898 172133 273134
rect 172369 272898 172425 273134
rect 172077 272866 172425 272898
rect 283921 273454 284269 273486
rect 283921 273218 283977 273454
rect 284213 273218 284269 273454
rect 283921 273134 284269 273218
rect 283921 272898 283977 273134
rect 284213 272898 284269 273134
rect 283921 272866 284269 272898
rect 378985 273454 379333 273486
rect 378985 273218 379041 273454
rect 379277 273218 379333 273454
rect 378985 273134 379333 273218
rect 378985 272898 379041 273134
rect 379277 272898 379333 273134
rect 378985 272866 379333 272898
rect 402468 273454 402868 273486
rect 402468 273218 402550 273454
rect 402786 273218 402868 273454
rect 402468 273134 402868 273218
rect 402468 272898 402550 273134
rect 402786 272898 402868 273134
rect 402468 272866 402868 272898
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 60412 255454 60812 255486
rect 60412 255218 60494 255454
rect 60730 255218 60812 255454
rect 60412 255134 60812 255218
rect 60412 254898 60494 255134
rect 60730 254898 60812 255134
rect 60412 254866 60812 254898
rect 77693 255454 78041 255486
rect 77693 255218 77749 255454
rect 77985 255218 78041 255454
rect 77693 255134 78041 255218
rect 77693 254898 77749 255134
rect 77985 254898 78041 255134
rect 77693 254866 78041 254898
rect 171397 255454 171745 255486
rect 171397 255218 171453 255454
rect 171689 255218 171745 255454
rect 171397 255134 171745 255218
rect 171397 254898 171453 255134
rect 171689 254898 171745 255134
rect 171397 254866 171745 254898
rect 284601 255454 284949 255486
rect 284601 255218 284657 255454
rect 284893 255218 284949 255454
rect 284601 255134 284949 255218
rect 284601 254898 284657 255134
rect 284893 254898 284949 255134
rect 284601 254866 284949 254898
rect 378305 255454 378653 255486
rect 378305 255218 378361 255454
rect 378597 255218 378653 255454
rect 378305 255134 378653 255218
rect 378305 254898 378361 255134
rect 378597 254898 378653 255134
rect 378305 254866 378653 254898
rect 403268 255454 403668 255486
rect 403268 255218 403350 255454
rect 403586 255218 403668 255454
rect 403268 255134 403668 255218
rect 403268 254898 403350 255134
rect 403586 254898 403668 255134
rect 403268 254866 403668 254898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 61212 237454 61612 237486
rect 61212 237218 61294 237454
rect 61530 237218 61612 237454
rect 61212 237134 61612 237218
rect 61212 236898 61294 237134
rect 61530 236898 61612 237134
rect 61212 236866 61612 236898
rect 77013 237454 77361 237486
rect 77013 237218 77069 237454
rect 77305 237218 77361 237454
rect 77013 237134 77361 237218
rect 77013 236898 77069 237134
rect 77305 236898 77361 237134
rect 77013 236866 77361 236898
rect 172077 237454 172425 237486
rect 172077 237218 172133 237454
rect 172369 237218 172425 237454
rect 172077 237134 172425 237218
rect 172077 236898 172133 237134
rect 172369 236898 172425 237134
rect 172077 236866 172425 236898
rect 283921 237454 284269 237486
rect 283921 237218 283977 237454
rect 284213 237218 284269 237454
rect 283921 237134 284269 237218
rect 283921 236898 283977 237134
rect 284213 236898 284269 237134
rect 283921 236866 284269 236898
rect 378985 237454 379333 237486
rect 378985 237218 379041 237454
rect 379277 237218 379333 237454
rect 378985 237134 379333 237218
rect 378985 236898 379041 237134
rect 379277 236898 379333 237134
rect 378985 236866 379333 236898
rect 402468 237454 402868 237486
rect 402468 237218 402550 237454
rect 402786 237218 402868 237454
rect 402468 237134 402868 237218
rect 402468 236898 402550 237134
rect 402786 236898 402868 237134
rect 402468 236866 402868 236898
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 60412 219454 60812 219486
rect 60412 219218 60494 219454
rect 60730 219218 60812 219454
rect 60412 219134 60812 219218
rect 60412 218898 60494 219134
rect 60730 218898 60812 219134
rect 60412 218866 60812 218898
rect 77693 219454 78041 219486
rect 77693 219218 77749 219454
rect 77985 219218 78041 219454
rect 77693 219134 78041 219218
rect 77693 218898 77749 219134
rect 77985 218898 78041 219134
rect 77693 218866 78041 218898
rect 171397 219454 171745 219486
rect 171397 219218 171453 219454
rect 171689 219218 171745 219454
rect 171397 219134 171745 219218
rect 171397 218898 171453 219134
rect 171689 218898 171745 219134
rect 171397 218866 171745 218898
rect 284601 219454 284949 219486
rect 284601 219218 284657 219454
rect 284893 219218 284949 219454
rect 284601 219134 284949 219218
rect 284601 218898 284657 219134
rect 284893 218898 284949 219134
rect 284601 218866 284949 218898
rect 378305 219454 378653 219486
rect 378305 219218 378361 219454
rect 378597 219218 378653 219454
rect 378305 219134 378653 219218
rect 378305 218898 378361 219134
rect 378597 218898 378653 219134
rect 378305 218866 378653 218898
rect 403268 219454 403668 219486
rect 403268 219218 403350 219454
rect 403586 219218 403668 219454
rect 403268 219134 403668 219218
rect 403268 218898 403350 219134
rect 403586 218898 403668 219134
rect 403268 218866 403668 218898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 61212 201454 61612 201486
rect 61212 201218 61294 201454
rect 61530 201218 61612 201454
rect 61212 201134 61612 201218
rect 61212 200898 61294 201134
rect 61530 200898 61612 201134
rect 61212 200866 61612 200898
rect 283921 201454 284269 201486
rect 283921 201218 283977 201454
rect 284213 201218 284269 201454
rect 283921 201134 284269 201218
rect 283921 200898 283977 201134
rect 284213 200898 284269 201134
rect 283921 200866 284269 200898
rect 378985 201454 379333 201486
rect 378985 201218 379041 201454
rect 379277 201218 379333 201454
rect 378985 201134 379333 201218
rect 378985 200898 379041 201134
rect 379277 200898 379333 201134
rect 378985 200866 379333 200898
rect 402468 201454 402868 201486
rect 402468 201218 402550 201454
rect 402786 201218 402868 201454
rect 402468 201134 402868 201218
rect 402468 200898 402550 201134
rect 402786 200898 402868 201134
rect 402468 200866 402868 200898
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 60412 183454 60812 183486
rect 60412 183218 60494 183454
rect 60730 183218 60812 183454
rect 60412 183134 60812 183218
rect 60412 182898 60494 183134
rect 60730 182898 60812 183134
rect 60412 182866 60812 182898
rect 403268 183454 403668 183486
rect 403268 183218 403350 183454
rect 403586 183218 403668 183454
rect 403268 183134 403668 183218
rect 403268 182898 403350 183134
rect 403586 182898 403668 183134
rect 403268 182866 403668 182898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 61212 165454 61612 165486
rect 61212 165218 61294 165454
rect 61530 165218 61612 165454
rect 61212 165134 61612 165218
rect 61212 164898 61294 165134
rect 61530 164898 61612 165134
rect 61212 164866 61612 164898
rect 402468 165454 402868 165486
rect 402468 165218 402550 165454
rect 402786 165218 402868 165454
rect 402468 165134 402868 165218
rect 402468 164898 402550 165134
rect 402786 164898 402868 165134
rect 402468 164866 402868 164898
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 60412 147454 60812 147486
rect 60412 147218 60494 147454
rect 60730 147218 60812 147454
rect 60412 147134 60812 147218
rect 60412 146898 60494 147134
rect 60730 146898 60812 147134
rect 60412 146866 60812 146898
rect 403268 147454 403668 147486
rect 403268 147218 403350 147454
rect 403586 147218 403668 147454
rect 403268 147134 403668 147218
rect 403268 146898 403350 147134
rect 403586 146898 403668 147134
rect 403268 146866 403668 146898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 61212 129454 61612 129486
rect 61212 129218 61294 129454
rect 61530 129218 61612 129454
rect 61212 129134 61612 129218
rect 61212 128898 61294 129134
rect 61530 128898 61612 129134
rect 61212 128866 61612 128898
rect 402468 129454 402868 129486
rect 402468 129218 402550 129454
rect 402786 129218 402868 129454
rect 402468 129134 402868 129218
rect 402468 128898 402550 129134
rect 402786 128898 402868 129134
rect 402468 128866 402868 128898
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 60412 111454 60812 111486
rect 60412 111218 60494 111454
rect 60730 111218 60812 111454
rect 60412 111134 60812 111218
rect 60412 110898 60494 111134
rect 60730 110898 60812 111134
rect 60412 110866 60812 110898
rect 403268 111454 403668 111486
rect 403268 111218 403350 111454
rect 403586 111218 403668 111454
rect 403268 111134 403668 111218
rect 403268 110898 403350 111134
rect 403586 110898 403668 111134
rect 403268 110866 403668 110898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 61212 93454 61612 93486
rect 61212 93218 61294 93454
rect 61530 93218 61612 93454
rect 61212 93134 61612 93218
rect 61212 92898 61294 93134
rect 61530 92898 61612 93134
rect 61212 92866 61612 92898
rect 402468 93454 402868 93486
rect 402468 93218 402550 93454
rect 402786 93218 402868 93454
rect 402468 93134 402868 93218
rect 402468 92898 402550 93134
rect 402786 92898 402868 93134
rect 402468 92866 402868 92898
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 60412 75454 60812 75486
rect 60412 75218 60494 75454
rect 60730 75218 60812 75454
rect 60412 75134 60812 75218
rect 60412 74898 60494 75134
rect 60730 74898 60812 75134
rect 60412 74866 60812 74898
rect 403268 75454 403668 75486
rect 403268 75218 403350 75454
rect 403586 75218 403668 75454
rect 403268 75134 403668 75218
rect 403268 74898 403350 75134
rect 403586 74898 403668 75134
rect 403268 74866 403668 74898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 61174 60134 70000
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 64894 63854 70000
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 70000
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 70000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 70000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 70000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 70000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 70000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 70000
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 70000
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 70000
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 70000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 70000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 70000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 70000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 70000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 70000
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 70000
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 70000
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 70000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 70000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 70000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 70000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 70000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 70000
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 70000
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 68614 175574 70000
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 70000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 70000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 70000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 70000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 70000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 61174 204134 70000
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 70000
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 70000
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 70000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 70000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 70000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 70000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 70000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 70000
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 70000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 70000
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 70000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 70000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 70000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 70000
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57454 272414 70000
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 70000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 70000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 70000
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 70000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 70000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 70000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 70000
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 70000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 61174 312134 70000
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 64894 315854 70000
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 68614 319574 70000
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 70000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 70000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 70000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 70000
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 70000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 61174 348134 70000
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 64894 351854 70000
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 68614 355574 70000
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 70000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 70000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 70000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 70000
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 57454 380414 70000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 61174 384134 70000
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 64894 387854 70000
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 68614 391574 70000
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 70000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 70000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 70000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 60494 363218 60730 363454
rect 60494 362898 60730 363134
rect 403350 363218 403586 363454
rect 403350 362898 403586 363134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 61294 345218 61530 345454
rect 61294 344898 61530 345134
rect 402550 345218 402786 345454
rect 402550 344898 402786 345134
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 60494 327218 60730 327454
rect 60494 326898 60730 327134
rect 403350 327218 403586 327454
rect 403350 326898 403586 327134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 61294 309218 61530 309454
rect 61294 308898 61530 309134
rect 402550 309218 402786 309454
rect 402550 308898 402786 309134
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 60494 291218 60730 291454
rect 60494 290898 60730 291134
rect 403350 291218 403586 291454
rect 403350 290898 403586 291134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 61294 273218 61530 273454
rect 61294 272898 61530 273134
rect 77069 273218 77305 273454
rect 77069 272898 77305 273134
rect 172133 273218 172369 273454
rect 172133 272898 172369 273134
rect 283977 273218 284213 273454
rect 283977 272898 284213 273134
rect 379041 273218 379277 273454
rect 379041 272898 379277 273134
rect 402550 273218 402786 273454
rect 402550 272898 402786 273134
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 60494 255218 60730 255454
rect 60494 254898 60730 255134
rect 77749 255218 77985 255454
rect 77749 254898 77985 255134
rect 171453 255218 171689 255454
rect 171453 254898 171689 255134
rect 284657 255218 284893 255454
rect 284657 254898 284893 255134
rect 378361 255218 378597 255454
rect 378361 254898 378597 255134
rect 403350 255218 403586 255454
rect 403350 254898 403586 255134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 61294 237218 61530 237454
rect 61294 236898 61530 237134
rect 77069 237218 77305 237454
rect 77069 236898 77305 237134
rect 172133 237218 172369 237454
rect 172133 236898 172369 237134
rect 283977 237218 284213 237454
rect 283977 236898 284213 237134
rect 379041 237218 379277 237454
rect 379041 236898 379277 237134
rect 402550 237218 402786 237454
rect 402550 236898 402786 237134
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 60494 219218 60730 219454
rect 60494 218898 60730 219134
rect 77749 219218 77985 219454
rect 77749 218898 77985 219134
rect 171453 219218 171689 219454
rect 171453 218898 171689 219134
rect 284657 219218 284893 219454
rect 284657 218898 284893 219134
rect 378361 219218 378597 219454
rect 378361 218898 378597 219134
rect 403350 219218 403586 219454
rect 403350 218898 403586 219134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 61294 201218 61530 201454
rect 61294 200898 61530 201134
rect 283977 201218 284213 201454
rect 283977 200898 284213 201134
rect 379041 201218 379277 201454
rect 379041 200898 379277 201134
rect 402550 201218 402786 201454
rect 402550 200898 402786 201134
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 60494 183218 60730 183454
rect 60494 182898 60730 183134
rect 403350 183218 403586 183454
rect 403350 182898 403586 183134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 61294 165218 61530 165454
rect 61294 164898 61530 165134
rect 402550 165218 402786 165454
rect 402550 164898 402786 165134
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 60494 147218 60730 147454
rect 60494 146898 60730 147134
rect 403350 147218 403586 147454
rect 403350 146898 403586 147134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 61294 129218 61530 129454
rect 61294 128898 61530 129134
rect 402550 129218 402786 129454
rect 402550 128898 402786 129134
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 60494 111218 60730 111454
rect 60494 110898 60730 111134
rect 403350 111218 403586 111454
rect 403350 110898 403586 111134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 61294 93218 61530 93454
rect 61294 92898 61530 93134
rect 402550 93218 402786 93454
rect 402550 92898 402786 93134
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 60494 75218 60730 75454
rect 60494 74898 60730 75134
rect 403350 75218 403586 75454
rect 403350 74898 403586 75134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 60494 363454
rect 60730 363218 403350 363454
rect 403586 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 60494 363134
rect 60730 362898 403350 363134
rect 403586 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 61294 345454
rect 61530 345218 402550 345454
rect 402786 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 61294 345134
rect 61530 344898 402550 345134
rect 402786 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 60494 327454
rect 60730 327218 403350 327454
rect 403586 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 60494 327134
rect 60730 326898 403350 327134
rect 403586 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 61294 309454
rect 61530 309218 402550 309454
rect 402786 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 61294 309134
rect 61530 308898 402550 309134
rect 402786 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 60494 291454
rect 60730 291218 403350 291454
rect 403586 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 60494 291134
rect 60730 290898 403350 291134
rect 403586 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 61294 273454
rect 61530 273218 77069 273454
rect 77305 273218 172133 273454
rect 172369 273218 283977 273454
rect 284213 273218 379041 273454
rect 379277 273218 402550 273454
rect 402786 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 61294 273134
rect 61530 272898 77069 273134
rect 77305 272898 172133 273134
rect 172369 272898 283977 273134
rect 284213 272898 379041 273134
rect 379277 272898 402550 273134
rect 402786 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 60494 255454
rect 60730 255218 77749 255454
rect 77985 255218 171453 255454
rect 171689 255218 284657 255454
rect 284893 255218 378361 255454
rect 378597 255218 403350 255454
rect 403586 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 60494 255134
rect 60730 254898 77749 255134
rect 77985 254898 171453 255134
rect 171689 254898 284657 255134
rect 284893 254898 378361 255134
rect 378597 254898 403350 255134
rect 403586 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 61294 237454
rect 61530 237218 77069 237454
rect 77305 237218 172133 237454
rect 172369 237218 283977 237454
rect 284213 237218 379041 237454
rect 379277 237218 402550 237454
rect 402786 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 61294 237134
rect 61530 236898 77069 237134
rect 77305 236898 172133 237134
rect 172369 236898 283977 237134
rect 284213 236898 379041 237134
rect 379277 236898 402550 237134
rect 402786 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 60494 219454
rect 60730 219218 77749 219454
rect 77985 219218 171453 219454
rect 171689 219218 284657 219454
rect 284893 219218 378361 219454
rect 378597 219218 403350 219454
rect 403586 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 60494 219134
rect 60730 218898 77749 219134
rect 77985 218898 171453 219134
rect 171689 218898 284657 219134
rect 284893 218898 378361 219134
rect 378597 218898 403350 219134
rect 403586 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 61294 201454
rect 61530 201218 283977 201454
rect 284213 201218 379041 201454
rect 379277 201218 402550 201454
rect 402786 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 61294 201134
rect 61530 200898 283977 201134
rect 284213 200898 379041 201134
rect 379277 200898 402550 201134
rect 402786 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 60494 183454
rect 60730 183218 403350 183454
rect 403586 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 60494 183134
rect 60730 182898 403350 183134
rect 403586 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 61294 165454
rect 61530 165218 402550 165454
rect 402786 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 61294 165134
rect 61530 164898 402550 165134
rect 402786 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 60494 147454
rect 60730 147218 403350 147454
rect 403586 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 60494 147134
rect 60730 146898 403350 147134
rect 403586 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 61294 129454
rect 61530 129218 402550 129454
rect 402786 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 61294 129134
rect 61530 128898 402550 129134
rect 402786 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 60494 111454
rect 60730 111218 403350 111454
rect 403586 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 60494 111134
rect 60730 110898 403350 111134
rect 403586 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 61294 93454
rect 61530 93218 402550 93454
rect 402786 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 61294 93134
rect 61530 92898 402550 93134
rect 402786 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 60494 75454
rect 60730 75218 403350 75454
rect 403586 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 60494 75134
rect 60730 74898 403350 75134
rect 403586 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use azadi_soc_top_caravel  mprj
<<<<<<< HEAD
timestamp 1640101730
=======
timestamp 1640019720
>>>>>>> 931d98e1c1894db8467f2b2099012c09581bc7c4
transform 1 0 60000 0 1 72000
box 0 0 344080 293964
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 70000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 70000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 70000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 70000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 70000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 70000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 70000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 70000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 70000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 70000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 367964 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 367964 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 367964 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 367964 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 367964 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 367964 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 367964 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 367964 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 367964 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 367964 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 70000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 70000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 70000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 70000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 70000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 70000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 70000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 70000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 70000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 70000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 367964 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 367964 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 367964 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 367964 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 367964 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 367964 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 367964 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 367964 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 367964 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 367964 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 70000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 70000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 70000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 70000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 70000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 70000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 70000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 70000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 70000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 70000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 367964 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 367964 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 367964 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 367964 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 367964 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 367964 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 367964 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 367964 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 367964 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 367964 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 70000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 70000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 70000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 70000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 70000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 70000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 70000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 70000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 70000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 367964 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 367964 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 367964 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 367964 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 367964 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 367964 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 367964 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 367964 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 367964 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 70000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 70000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 70000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 70000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 70000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 70000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 70000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 70000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 70000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 70000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 367964 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 367964 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 367964 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 367964 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 367964 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 367964 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 367964 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 367964 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 367964 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 367964 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 70000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 70000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 70000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 70000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 70000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 70000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 70000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 70000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 70000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 70000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 367964 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 367964 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 367964 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 367964 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 367964 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 367964 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 367964 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 367964 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 367964 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 367964 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 70000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 70000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 70000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 70000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 70000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 70000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 70000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 70000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 70000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 367964 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 367964 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 367964 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 367964 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 367964 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 367964 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 367964 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 367964 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 367964 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 70000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 70000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 70000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 70000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 70000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 70000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 70000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 70000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 70000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 70000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 367964 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 367964 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 367964 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 367964 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 367964 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 367964 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 367964 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 367964 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 367964 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 367964 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
