##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Fri Dec 17 18:10:46 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 1720.400000 BY 1469.820000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.420000 0.000000 3.560000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.540000 0.000000 1.680000 0.490000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.785000 0.000000 362.925000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.045000 0.000000 122.185000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.275000 0.000000 366.415000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.295000 0.000000 359.435000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.810000 0.000000 355.950000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.320000 0.000000 352.460000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.830000 0.000000 348.970000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.695000 0.000000 233.835000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.205000 0.000000 230.345000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.715000 0.000000 226.855000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.225000 0.000000 223.365000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.735000 0.000000 219.875000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.250000 0.000000 216.390000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.760000 0.000000 212.900000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.270000 0.000000 209.410000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.780000 0.000000 205.920000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.290000 0.000000 202.430000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.805000 0.000000 198.945000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.315000 0.000000 195.455000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.825000 0.000000 191.965000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.335000 0.000000 188.475000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.845000 0.000000 184.985000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.360000 0.000000 181.500000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.870000 0.000000 178.010000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.380000 0.000000 174.520000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.890000 0.000000 171.030000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.400000 0.000000 167.540000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.915000 0.000000 164.055000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.425000 0.000000 160.565000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.935000 0.000000 157.075000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.445000 0.000000 153.585000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.955000 0.000000 150.095000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.470000 0.000000 146.610000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.980000 0.000000 143.120000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.490000 0.000000 139.630000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.000000 0.000000 136.140000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.510000 0.000000 132.650000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.025000 0.000000 129.165000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.535000 0.000000 125.675000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.555000 0.000000 118.695000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.065000 0.000000 115.205000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.580000 0.000000 111.720000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.090000 0.000000 108.230000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.600000 0.000000 104.740000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.110000 0.000000 101.250000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.620000 0.000000 97.760000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.135000 0.000000 94.275000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.645000 0.000000 90.785000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.155000 0.000000 87.295000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.665000 0.000000 83.805000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.175000 0.000000 80.315000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.690000 0.000000 76.830000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.200000 0.000000 73.340000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.710000 0.000000 69.850000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.220000 0.000000 66.360000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.730000 0.000000 62.870000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.245000 0.000000 59.385000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.755000 0.000000 55.895000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.265000 0.000000 52.405000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.775000 0.000000 48.915000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.285000 0.000000 45.425000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.800000 0.000000 41.940000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.310000 0.000000 38.450000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.820000 0.000000 34.960000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.330000 0.000000 31.470000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.840000 0.000000 27.980000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.355000 0.000000 24.495000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.865000 0.000000 21.005000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.375000 0.000000 17.515000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.885000 0.000000 14.025000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.395000 0.000000 10.535000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.910000 0.000000 7.050000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.340000 0.000000 345.480000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.850000 0.000000 341.990000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.365000 0.000000 338.505000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.875000 0.000000 335.015000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.385000 0.000000 331.525000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.895000 0.000000 328.035000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.405000 0.000000 324.545000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.920000 0.000000 321.060000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.430000 0.000000 317.570000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.940000 0.000000 314.080000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.450000 0.000000 310.590000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.960000 0.000000 307.100000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.475000 0.000000 303.615000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.985000 0.000000 300.125000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.495000 0.000000 296.635000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.005000 0.000000 293.145000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.515000 0.000000 289.655000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.030000 0.000000 286.170000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.540000 0.000000 282.680000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.050000 0.000000 279.190000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.560000 0.000000 275.700000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.070000 0.000000 272.210000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.585000 0.000000 268.725000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.095000 0.000000 265.235000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.605000 0.000000 261.745000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.115000 0.000000 258.255000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.625000 0.000000 254.765000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.140000 0.000000 251.280000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.650000 0.000000 247.790000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.160000 0.000000 244.300000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670000 0.000000 240.810000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.180000 0.000000 237.320000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.865000 0.000000 813.005000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.380000 0.000000 809.520000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.890000 0.000000 806.030000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.400000 0.000000 802.540000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.910000 0.000000 799.050000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.420000 0.000000 795.560000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.935000 0.000000 792.075000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.445000 0.000000 788.585000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.955000 0.000000 785.095000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.465000 0.000000 781.605000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.975000 0.000000 778.115000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.490000 0.000000 774.630000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.000000 0.000000 771.140000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.510000 0.000000 767.650000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.020000 0.000000 764.160000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.530000 0.000000 760.670000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.045000 0.000000 757.185000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.555000 0.000000 753.695000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.065000 0.000000 750.205000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.575000 0.000000 746.715000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.085000 0.000000 743.225000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.600000 0.000000 739.740000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.110000 0.000000 736.250000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.620000 0.000000 732.760000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.130000 0.000000 729.270000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.640000 0.000000 725.780000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.155000 0.000000 722.295000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.665000 0.000000 718.805000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.175000 0.000000 715.315000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.685000 0.000000 711.825000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.195000 0.000000 708.335000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.710000 0.000000 704.850000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.220000 0.000000 701.360000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.730000 0.000000 697.870000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.240000 0.000000 694.380000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.750000 0.000000 690.890000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.265000 0.000000 687.405000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.775000 0.000000 683.915000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.285000 0.000000 680.425000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.795000 0.000000 676.935000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.305000 0.000000 673.445000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.820000 0.000000 669.960000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.330000 0.000000 666.470000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.840000 0.000000 662.980000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.350000 0.000000 659.490000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.860000 0.000000 656.000000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.375000 0.000000 652.515000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.885000 0.000000 649.025000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.395000 0.000000 645.535000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.905000 0.000000 642.045000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.415000 0.000000 638.555000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.930000 0.000000 635.070000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.440000 0.000000 631.580000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.950000 0.000000 628.090000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.460000 0.000000 624.600000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.970000 0.000000 621.110000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.485000 0.000000 617.625000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.995000 0.000000 614.135000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.505000 0.000000 610.645000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.015000 0.000000 607.155000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.525000 0.000000 603.665000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.040000 0.000000 600.180000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.550000 0.000000 596.690000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.060000 0.000000 593.200000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.570000 0.000000 589.710000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.080000 0.000000 586.220000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.595000 0.000000 582.735000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.105000 0.000000 579.245000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.615000 0.000000 575.755000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.125000 0.000000 572.265000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.635000 0.000000 568.775000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.150000 0.000000 565.290000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.660000 0.000000 561.800000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.170000 0.000000 558.310000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.680000 0.000000 554.820000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.190000 0.000000 551.330000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.705000 0.000000 547.845000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.215000 0.000000 544.355000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.725000 0.000000 540.865000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.235000 0.000000 537.375000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.745000 0.000000 533.885000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.260000 0.000000 530.400000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.770000 0.000000 526.910000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.280000 0.000000 523.420000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.790000 0.000000 519.930000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.300000 0.000000 516.440000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.815000 0.000000 512.955000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.325000 0.000000 509.465000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.835000 0.000000 505.975000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.345000 0.000000 502.485000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.855000 0.000000 498.995000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.370000 0.000000 495.510000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.880000 0.000000 492.020000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.390000 0.000000 488.530000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.900000 0.000000 485.040000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.410000 0.000000 481.550000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.925000 0.000000 478.065000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.435000 0.000000 474.575000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.945000 0.000000 471.085000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.455000 0.000000 467.595000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.965000 0.000000 464.105000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.480000 0.000000 460.620000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.990000 0.000000 457.130000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.500000 0.000000 453.640000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.010000 0.000000 450.150000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.520000 0.000000 446.660000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.035000 0.000000 443.175000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.545000 0.000000 439.685000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.055000 0.000000 436.195000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.565000 0.000000 432.705000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.075000 0.000000 429.215000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590000 0.000000 425.730000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.100000 0.000000 422.240000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.610000 0.000000 418.750000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.120000 0.000000 415.260000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.630000 0.000000 411.770000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.145000 0.000000 408.285000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.655000 0.000000 404.795000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.165000 0.000000 401.305000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.675000 0.000000 397.815000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.185000 0.000000 394.325000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.700000 0.000000 390.840000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.210000 0.000000 387.350000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.720000 0.000000 383.860000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.230000 0.000000 380.370000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.740000 0.000000 376.880000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.255000 0.000000 373.395000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.765000 0.000000 369.905000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.460000 0.000000 1259.600000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.970000 0.000000 1256.110000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.480000 0.000000 1252.620000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.990000 0.000000 1249.130000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.505000 0.000000 1245.645000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.015000 0.000000 1242.155000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.525000 0.000000 1238.665000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.035000 0.000000 1235.175000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.545000 0.000000 1231.685000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.060000 0.000000 1228.200000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.570000 0.000000 1224.710000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.080000 0.000000 1221.220000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.590000 0.000000 1217.730000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.100000 0.000000 1214.240000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.615000 0.000000 1210.755000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.125000 0.000000 1207.265000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.635000 0.000000 1203.775000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.145000 0.000000 1200.285000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.655000 0.000000 1196.795000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.170000 0.000000 1193.310000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.680000 0.000000 1189.820000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.190000 0.000000 1186.330000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.700000 0.000000 1182.840000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.210000 0.000000 1179.350000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.725000 0.000000 1175.865000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.235000 0.000000 1172.375000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.745000 0.000000 1168.885000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.255000 0.000000 1165.395000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.765000 0.000000 1161.905000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.280000 0.000000 1158.420000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.790000 0.000000 1154.930000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.300000 0.000000 1151.440000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.810000 0.000000 1147.950000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.320000 0.000000 1144.460000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.835000 0.000000 1140.975000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.345000 0.000000 1137.485000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.855000 0.000000 1133.995000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.365000 0.000000 1130.505000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.875000 0.000000 1127.015000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.390000 0.000000 1123.530000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.900000 0.000000 1120.040000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.410000 0.000000 1116.550000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.920000 0.000000 1113.060000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.430000 0.000000 1109.570000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.945000 0.000000 1106.085000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.455000 0.000000 1102.595000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.965000 0.000000 1099.105000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.475000 0.000000 1095.615000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.985000 0.000000 1092.125000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.500000 0.000000 1088.640000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.010000 0.000000 1085.150000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.520000 0.000000 1081.660000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.030000 0.000000 1078.170000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.540000 0.000000 1074.680000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.055000 0.000000 1071.195000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.565000 0.000000 1067.705000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.075000 0.000000 1064.215000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.585000 0.000000 1060.725000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.095000 0.000000 1057.235000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.610000 0.000000 1053.750000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.120000 0.000000 1050.260000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.630000 0.000000 1046.770000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.140000 0.000000 1043.280000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.650000 0.000000 1039.790000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.165000 0.000000 1036.305000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.675000 0.000000 1032.815000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.185000 0.000000 1029.325000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.695000 0.000000 1025.835000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.205000 0.000000 1022.345000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.720000 0.000000 1018.860000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.230000 0.000000 1015.370000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.740000 0.000000 1011.880000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.250000 0.000000 1008.390000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.760000 0.000000 1004.900000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.275000 0.000000 1001.415000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.785000 0.000000 997.925000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.295000 0.000000 994.435000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.805000 0.000000 990.945000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.315000 0.000000 987.455000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.830000 0.000000 983.970000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.340000 0.000000 980.480000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.850000 0.000000 976.990000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.360000 0.000000 973.500000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.870000 0.000000 970.010000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.385000 0.000000 966.525000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.895000 0.000000 963.035000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.405000 0.000000 959.545000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.915000 0.000000 956.055000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.425000 0.000000 952.565000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.940000 0.000000 949.080000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.450000 0.000000 945.590000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.960000 0.000000 942.100000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.470000 0.000000 938.610000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.980000 0.000000 935.120000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.495000 0.000000 931.635000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.005000 0.000000 928.145000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.515000 0.000000 924.655000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.025000 0.000000 921.165000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.535000 0.000000 917.675000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.050000 0.000000 914.190000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.560000 0.000000 910.700000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070000 0.000000 907.210000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.580000 0.000000 903.720000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.090000 0.000000 900.230000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.605000 0.000000 896.745000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.115000 0.000000 893.255000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.625000 0.000000 889.765000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.135000 0.000000 886.275000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.645000 0.000000 882.785000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.160000 0.000000 879.300000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.670000 0.000000 875.810000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.180000 0.000000 872.320000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.690000 0.000000 868.830000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.200000 0.000000 865.340000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.715000 0.000000 861.855000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.225000 0.000000 858.365000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.735000 0.000000 854.875000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.245000 0.000000 851.385000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.755000 0.000000 847.895000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.270000 0.000000 844.410000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.780000 0.000000 840.920000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290000 0.000000 837.430000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.800000 0.000000 833.940000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.310000 0.000000 830.450000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.825000 0.000000 826.965000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.335000 0.000000 823.475000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.845000 0.000000 819.985000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.355000 0.000000 816.495000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.050000 0.000000 1706.190000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.560000 0.000000 1702.700000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.075000 0.000000 1699.215000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1695.585000 0.000000 1695.725000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.095000 0.000000 1692.235000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.605000 0.000000 1688.745000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.115000 0.000000 1685.255000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.630000 0.000000 1681.770000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.140000 0.000000 1678.280000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.650000 0.000000 1674.790000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.160000 0.000000 1671.300000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.670000 0.000000 1667.810000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.185000 0.000000 1664.325000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.695000 0.000000 1660.835000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.205000 0.000000 1657.345000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.715000 0.000000 1653.855000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.225000 0.000000 1650.365000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.740000 0.000000 1646.880000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.250000 0.000000 1643.390000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.760000 0.000000 1639.900000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.270000 0.000000 1636.410000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.780000 0.000000 1632.920000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.295000 0.000000 1629.435000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.805000 0.000000 1625.945000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.315000 0.000000 1622.455000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.825000 0.000000 1618.965000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.335000 0.000000 1615.475000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.850000 0.000000 1611.990000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1608.360000 0.000000 1608.500000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.870000 0.000000 1605.010000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1601.380000 0.000000 1601.520000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.890000 0.000000 1598.030000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.405000 0.000000 1594.545000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.915000 0.000000 1591.055000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.425000 0.000000 1587.565000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.935000 0.000000 1584.075000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.445000 0.000000 1580.585000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.960000 0.000000 1577.100000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.470000 0.000000 1573.610000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.980000 0.000000 1570.120000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.490000 0.000000 1566.630000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.000000 0.000000 1563.140000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.515000 0.000000 1559.655000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.025000 0.000000 1556.165000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.535000 0.000000 1552.675000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.045000 0.000000 1549.185000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.555000 0.000000 1545.695000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.070000 0.000000 1542.210000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.580000 0.000000 1538.720000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.090000 0.000000 1535.230000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.600000 0.000000 1531.740000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.110000 0.000000 1528.250000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.625000 0.000000 1524.765000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.135000 0.000000 1521.275000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.645000 0.000000 1517.785000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.155000 0.000000 1514.295000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.665000 0.000000 1510.805000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.180000 0.000000 1507.320000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690000 0.000000 1503.830000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.200000 0.000000 1500.340000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.710000 0.000000 1496.850000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.220000 0.000000 1493.360000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.735000 0.000000 1489.875000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.245000 0.000000 1486.385000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.755000 0.000000 1482.895000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.265000 0.000000 1479.405000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.775000 0.000000 1475.915000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.290000 0.000000 1472.430000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.800000 0.000000 1468.940000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.310000 0.000000 1465.450000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.820000 0.000000 1461.960000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.330000 0.000000 1458.470000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.845000 0.000000 1454.985000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.355000 0.000000 1451.495000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.865000 0.000000 1448.005000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.375000 0.000000 1444.515000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.885000 0.000000 1441.025000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.400000 0.000000 1437.540000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.910000 0.000000 1434.050000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1430.420000 0.000000 1430.560000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.930000 0.000000 1427.070000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.440000 0.000000 1423.580000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.955000 0.000000 1420.095000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.465000 0.000000 1416.605000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.975000 0.000000 1413.115000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.485000 0.000000 1409.625000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.995000 0.000000 1406.135000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.510000 0.000000 1402.650000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.020000 0.000000 1399.160000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.530000 0.000000 1395.670000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.040000 0.000000 1392.180000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.550000 0.000000 1388.690000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.065000 0.000000 1385.205000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.575000 0.000000 1381.715000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.085000 0.000000 1378.225000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.595000 0.000000 1374.735000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.105000 0.000000 1371.245000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.620000 0.000000 1367.760000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.130000 0.000000 1364.270000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.640000 0.000000 1360.780000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.150000 0.000000 1357.290000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.660000 0.000000 1353.800000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.175000 0.000000 1350.315000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.685000 0.000000 1346.825000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1343.195000 0.000000 1343.335000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.705000 0.000000 1339.845000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.215000 0.000000 1336.355000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.730000 0.000000 1332.870000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.240000 0.000000 1329.380000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.750000 0.000000 1325.890000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.260000 0.000000 1322.400000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.770000 0.000000 1318.910000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.285000 0.000000 1315.425000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.795000 0.000000 1311.935000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.305000 0.000000 1308.445000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.815000 0.000000 1304.955000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.325000 0.000000 1301.465000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.840000 0.000000 1297.980000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.350000 0.000000 1294.490000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.860000 0.000000 1291.000000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.370000 0.000000 1287.510000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.880000 0.000000 1284.020000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.395000 0.000000 1280.535000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.905000 0.000000 1277.045000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.415000 0.000000 1273.555000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.925000 0.000000 1270.065000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.435000 0.000000 1266.575000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.950000 0.000000 1263.090000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 55.315000 0.800000 55.615000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.510000 0.800000 138.810000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 221.705000 0.800000 222.005000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 332.635000 0.800000 332.935000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 443.560000 0.800000 443.860000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 554.490000 0.800000 554.790000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 665.420000 0.800000 665.720000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 776.345000 0.800000 776.645000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 887.275000 0.800000 887.575000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 998.200000 0.800000 998.500000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1109.130000 0.800000 1109.430000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1220.060000 0.800000 1220.360000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1330.985000 0.800000 1331.285000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1441.915000 0.800000 1442.215000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.390000 1469.330000 147.530000 1469.820000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.010000 1469.330000 344.150000 1469.820000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.625000 1469.330000 540.765000 1469.820000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.240000 1469.330000 737.380000 1469.820000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.855000 1469.330000 933.995000 1469.820000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.470000 1469.330000 1130.610000 1469.820000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.090000 1469.330000 1327.230000 1469.820000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.705000 1469.330000 1523.845000 1469.820000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.040000 1469.330000 1715.180000 1469.820000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1413.100000 1720.400000 1413.400000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1300.040000 1720.400000 1300.340000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1186.980000 1720.400000 1187.280000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1073.920000 1720.400000 1074.220000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 960.860000 1720.400000 961.160000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 847.800000 1720.400000 848.100000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 734.740000 1720.400000 735.040000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 621.680000 1720.400000 621.980000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 508.620000 1720.400000 508.920000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 423.825000 1720.400000 424.125000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 339.030000 1720.400000 339.330000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 254.235000 1720.400000 254.535000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 169.440000 1720.400000 169.740000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 84.645000 1720.400000 84.945000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 3.780000 1720.400000 4.080000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 27.580000 0.800000 27.880000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 110.780000 0.800000 111.080000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 193.975000 0.800000 194.275000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 304.900000 0.800000 305.200000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 415.830000 0.800000 416.130000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 526.760000 0.800000 527.060000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 637.685000 0.800000 637.985000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 748.615000 0.800000 748.915000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 859.540000 0.800000 859.840000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 970.470000 0.800000 970.770000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1081.400000 0.800000 1081.700000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1192.325000 0.800000 1192.625000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1303.255000 0.800000 1303.555000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1414.180000 0.800000 1414.480000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.240000 1469.330000 98.380000 1469.820000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.855000 1469.330000 294.995000 1469.820000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.470000 1469.330000 491.610000 1469.820000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.085000 1469.330000 688.225000 1469.820000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.700000 1469.330000 884.840000 1469.820000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.320000 1469.330000 1081.460000 1469.820000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.935000 1469.330000 1278.075000 1469.820000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.550000 1469.330000 1474.690000 1469.820000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.165000 1469.330000 1671.305000 1469.820000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1441.365000 1720.400000 1441.665000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1328.305000 1720.400000 1328.605000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1215.245000 1720.400000 1215.545000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1102.185000 1720.400000 1102.485000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 989.125000 1720.400000 989.425000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 876.065000 1720.400000 876.365000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 763.005000 1720.400000 763.305000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 649.945000 1720.400000 650.245000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 536.885000 1720.400000 537.185000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 452.090000 1720.400000 452.390000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 367.295000 1720.400000 367.595000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 282.500000 1720.400000 282.800000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 197.705000 1720.400000 198.005000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 112.910000 1720.400000 113.210000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 28.115000 1720.400000 28.415000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 4.390000 0.800000 4.690000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 83.045000 0.800000 83.345000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 166.240000 0.800000 166.540000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 277.170000 0.800000 277.470000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 388.100000 0.800000 388.400000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 499.025000 0.800000 499.325000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 609.955000 0.800000 610.255000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 720.880000 0.800000 721.180000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 831.810000 0.800000 832.110000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 942.740000 0.800000 943.040000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1053.665000 0.800000 1053.965000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1164.595000 0.800000 1164.895000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1275.520000 0.800000 1275.820000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1386.450000 0.800000 1386.750000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.085000 1469.330000 49.225000 1469.820000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.700000 1469.330000 245.840000 1469.820000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.315000 1469.330000 442.455000 1469.820000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.930000 1469.330000 639.070000 1469.820000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.550000 1469.330000 835.690000 1469.820000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.165000 1469.330000 1032.305000 1469.820000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.780000 1469.330000 1228.920000 1469.820000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.395000 1469.330000 1425.535000 1469.820000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.010000 1469.330000 1622.150000 1469.820000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1464.730000 1720.400000 1465.030000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1356.570000 1720.400000 1356.870000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1243.510000 1720.400000 1243.810000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1130.450000 1720.400000 1130.750000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1017.390000 1720.400000 1017.690000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 904.330000 1720.400000 904.630000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 791.270000 1720.400000 791.570000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 678.210000 1720.400000 678.510000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 565.150000 1720.400000 565.450000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 480.355000 1720.400000 480.655000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 395.560000 1720.400000 395.860000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 310.765000 1720.400000 311.065000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 225.970000 1720.400000 226.270000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 141.175000 1720.400000 141.475000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 56.380000 1720.400000 56.680000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 249.440000 0.800000 249.740000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 360.365000 0.800000 360.665000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 471.295000 0.800000 471.595000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 582.220000 0.800000 582.520000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 693.150000 0.800000 693.450000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 804.080000 0.800000 804.380000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 915.005000 0.800000 915.305000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1025.935000 0.800000 1026.235000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1136.860000 0.800000 1137.160000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1247.790000 0.800000 1248.090000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1358.720000 0.800000 1359.020000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1465.340000 0.800000 1465.640000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.545000 1469.330000 196.685000 1469.820000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.160000 1469.330000 393.300000 1469.820000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.780000 1469.330000 589.920000 1469.820000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.395000 1469.330000 786.535000 1469.820000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.010000 1469.330000 983.150000 1469.820000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.625000 1469.330000 1179.765000 1469.820000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.240000 1469.330000 1376.380000 1469.820000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.860000 1469.330000 1573.000000 1469.820000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.300000 1469.330000 4.440000 1469.820000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1384.835000 1720.400000 1385.135000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1271.775000 1720.400000 1272.075000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1158.715000 1720.400000 1159.015000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 1045.655000 1720.400000 1045.955000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 932.595000 1720.400000 932.895000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 819.535000 1720.400000 819.835000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 706.475000 1720.400000 706.775000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1719.600000 593.415000 1720.400000 593.715000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.540000 0.000000 1709.680000 0.490000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.580000 0.000000 1714.720000 0.490000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.520000 0.000000 1716.660000 0.490000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.030000 0.000000 1713.170000 0.490000 ;
    END
  END user_irq[0]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1716.340000 1.930000 1718.340000 1467.720000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.060000 1.930000 4.060000 1467.720000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1123.005000 632.850000 1124.745000 1020.830000 ;
      LAYER met4 ;
        RECT 1591.525000 632.850000 1593.265000 1020.830000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 556.985000 648.195000 558.725000 1036.175000 ;
      LAYER met4 ;
        RECT 88.465000 648.195000 90.205000 1036.175000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1712.340000 5.930000 1714.340000 1463.720000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.060000 5.930000 8.060000 1463.720000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1594.925000 629.450000 1596.665000 1024.230000 ;
      LAYER met4 ;
        RECT 1119.605000 629.450000 1121.345000 1024.230000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 85.065000 644.795000 86.805000 1039.575000 ;
      LAYER met4 ;
        RECT 560.385000 644.795000 562.125000 1039.575000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END VGND
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1720.400000 1469.820000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1720.400000 1469.820000 ;
    LAYER met2 ;
      RECT 1715.320000 1469.190000 1720.400000 1469.820000 ;
      RECT 1671.445000 1469.190000 1714.900000 1469.820000 ;
      RECT 1622.290000 1469.190000 1671.025000 1469.820000 ;
      RECT 1573.140000 1469.190000 1621.870000 1469.820000 ;
      RECT 1523.985000 1469.190000 1572.720000 1469.820000 ;
      RECT 1474.830000 1469.190000 1523.565000 1469.820000 ;
      RECT 1425.675000 1469.190000 1474.410000 1469.820000 ;
      RECT 1376.520000 1469.190000 1425.255000 1469.820000 ;
      RECT 1327.370000 1469.190000 1376.100000 1469.820000 ;
      RECT 1278.215000 1469.190000 1326.950000 1469.820000 ;
      RECT 1229.060000 1469.190000 1277.795000 1469.820000 ;
      RECT 1179.905000 1469.190000 1228.640000 1469.820000 ;
      RECT 1130.750000 1469.190000 1179.485000 1469.820000 ;
      RECT 1081.600000 1469.190000 1130.330000 1469.820000 ;
      RECT 1032.445000 1469.190000 1081.180000 1469.820000 ;
      RECT 983.290000 1469.190000 1032.025000 1469.820000 ;
      RECT 934.135000 1469.190000 982.870000 1469.820000 ;
      RECT 884.980000 1469.190000 933.715000 1469.820000 ;
      RECT 835.830000 1469.190000 884.560000 1469.820000 ;
      RECT 786.675000 1469.190000 835.410000 1469.820000 ;
      RECT 737.520000 1469.190000 786.255000 1469.820000 ;
      RECT 688.365000 1469.190000 737.100000 1469.820000 ;
      RECT 639.210000 1469.190000 687.945000 1469.820000 ;
      RECT 590.060000 1469.190000 638.790000 1469.820000 ;
      RECT 540.905000 1469.190000 589.640000 1469.820000 ;
      RECT 491.750000 1469.190000 540.485000 1469.820000 ;
      RECT 442.595000 1469.190000 491.330000 1469.820000 ;
      RECT 393.440000 1469.190000 442.175000 1469.820000 ;
      RECT 344.290000 1469.190000 393.020000 1469.820000 ;
      RECT 295.135000 1469.190000 343.870000 1469.820000 ;
      RECT 245.980000 1469.190000 294.715000 1469.820000 ;
      RECT 196.825000 1469.190000 245.560000 1469.820000 ;
      RECT 147.670000 1469.190000 196.405000 1469.820000 ;
      RECT 98.520000 1469.190000 147.250000 1469.820000 ;
      RECT 49.365000 1469.190000 98.100000 1469.820000 ;
      RECT 4.580000 1469.190000 48.945000 1469.820000 ;
      RECT 0.000000 1469.190000 4.160000 1469.820000 ;
      RECT 0.000000 0.630000 1720.400000 1469.190000 ;
      RECT 1716.800000 0.000000 1720.400000 0.630000 ;
      RECT 1714.860000 0.000000 1716.380000 0.630000 ;
      RECT 1713.310000 0.000000 1714.440000 0.630000 ;
      RECT 1709.820000 0.000000 1712.890000 0.630000 ;
      RECT 1706.330000 0.000000 1709.400000 0.630000 ;
      RECT 1702.840000 0.000000 1705.910000 0.630000 ;
      RECT 1699.355000 0.000000 1702.420000 0.630000 ;
      RECT 1695.865000 0.000000 1698.935000 0.630000 ;
      RECT 1692.375000 0.000000 1695.445000 0.630000 ;
      RECT 1688.885000 0.000000 1691.955000 0.630000 ;
      RECT 1685.395000 0.000000 1688.465000 0.630000 ;
      RECT 1681.910000 0.000000 1684.975000 0.630000 ;
      RECT 1678.420000 0.000000 1681.490000 0.630000 ;
      RECT 1674.930000 0.000000 1678.000000 0.630000 ;
      RECT 1671.440000 0.000000 1674.510000 0.630000 ;
      RECT 1667.950000 0.000000 1671.020000 0.630000 ;
      RECT 1664.465000 0.000000 1667.530000 0.630000 ;
      RECT 1660.975000 0.000000 1664.045000 0.630000 ;
      RECT 1657.485000 0.000000 1660.555000 0.630000 ;
      RECT 1653.995000 0.000000 1657.065000 0.630000 ;
      RECT 1650.505000 0.000000 1653.575000 0.630000 ;
      RECT 1647.020000 0.000000 1650.085000 0.630000 ;
      RECT 1643.530000 0.000000 1646.600000 0.630000 ;
      RECT 1640.040000 0.000000 1643.110000 0.630000 ;
      RECT 1636.550000 0.000000 1639.620000 0.630000 ;
      RECT 1633.060000 0.000000 1636.130000 0.630000 ;
      RECT 1629.575000 0.000000 1632.640000 0.630000 ;
      RECT 1626.085000 0.000000 1629.155000 0.630000 ;
      RECT 1622.595000 0.000000 1625.665000 0.630000 ;
      RECT 1619.105000 0.000000 1622.175000 0.630000 ;
      RECT 1615.615000 0.000000 1618.685000 0.630000 ;
      RECT 1612.130000 0.000000 1615.195000 0.630000 ;
      RECT 1608.640000 0.000000 1611.710000 0.630000 ;
      RECT 1605.150000 0.000000 1608.220000 0.630000 ;
      RECT 1601.660000 0.000000 1604.730000 0.630000 ;
      RECT 1598.170000 0.000000 1601.240000 0.630000 ;
      RECT 1594.685000 0.000000 1597.750000 0.630000 ;
      RECT 1591.195000 0.000000 1594.265000 0.630000 ;
      RECT 1587.705000 0.000000 1590.775000 0.630000 ;
      RECT 1584.215000 0.000000 1587.285000 0.630000 ;
      RECT 1580.725000 0.000000 1583.795000 0.630000 ;
      RECT 1577.240000 0.000000 1580.305000 0.630000 ;
      RECT 1573.750000 0.000000 1576.820000 0.630000 ;
      RECT 1570.260000 0.000000 1573.330000 0.630000 ;
      RECT 1566.770000 0.000000 1569.840000 0.630000 ;
      RECT 1563.280000 0.000000 1566.350000 0.630000 ;
      RECT 1559.795000 0.000000 1562.860000 0.630000 ;
      RECT 1556.305000 0.000000 1559.375000 0.630000 ;
      RECT 1552.815000 0.000000 1555.885000 0.630000 ;
      RECT 1549.325000 0.000000 1552.395000 0.630000 ;
      RECT 1545.835000 0.000000 1548.905000 0.630000 ;
      RECT 1542.350000 0.000000 1545.415000 0.630000 ;
      RECT 1538.860000 0.000000 1541.930000 0.630000 ;
      RECT 1535.370000 0.000000 1538.440000 0.630000 ;
      RECT 1531.880000 0.000000 1534.950000 0.630000 ;
      RECT 1528.390000 0.000000 1531.460000 0.630000 ;
      RECT 1524.905000 0.000000 1527.970000 0.630000 ;
      RECT 1521.415000 0.000000 1524.485000 0.630000 ;
      RECT 1517.925000 0.000000 1520.995000 0.630000 ;
      RECT 1514.435000 0.000000 1517.505000 0.630000 ;
      RECT 1510.945000 0.000000 1514.015000 0.630000 ;
      RECT 1507.460000 0.000000 1510.525000 0.630000 ;
      RECT 1503.970000 0.000000 1507.040000 0.630000 ;
      RECT 1500.480000 0.000000 1503.550000 0.630000 ;
      RECT 1496.990000 0.000000 1500.060000 0.630000 ;
      RECT 1493.500000 0.000000 1496.570000 0.630000 ;
      RECT 1490.015000 0.000000 1493.080000 0.630000 ;
      RECT 1486.525000 0.000000 1489.595000 0.630000 ;
      RECT 1483.035000 0.000000 1486.105000 0.630000 ;
      RECT 1479.545000 0.000000 1482.615000 0.630000 ;
      RECT 1476.055000 0.000000 1479.125000 0.630000 ;
      RECT 1472.570000 0.000000 1475.635000 0.630000 ;
      RECT 1469.080000 0.000000 1472.150000 0.630000 ;
      RECT 1465.590000 0.000000 1468.660000 0.630000 ;
      RECT 1462.100000 0.000000 1465.170000 0.630000 ;
      RECT 1458.610000 0.000000 1461.680000 0.630000 ;
      RECT 1455.125000 0.000000 1458.190000 0.630000 ;
      RECT 1451.635000 0.000000 1454.705000 0.630000 ;
      RECT 1448.145000 0.000000 1451.215000 0.630000 ;
      RECT 1444.655000 0.000000 1447.725000 0.630000 ;
      RECT 1441.165000 0.000000 1444.235000 0.630000 ;
      RECT 1437.680000 0.000000 1440.745000 0.630000 ;
      RECT 1434.190000 0.000000 1437.260000 0.630000 ;
      RECT 1430.700000 0.000000 1433.770000 0.630000 ;
      RECT 1427.210000 0.000000 1430.280000 0.630000 ;
      RECT 1423.720000 0.000000 1426.790000 0.630000 ;
      RECT 1420.235000 0.000000 1423.300000 0.630000 ;
      RECT 1416.745000 0.000000 1419.815000 0.630000 ;
      RECT 1413.255000 0.000000 1416.325000 0.630000 ;
      RECT 1409.765000 0.000000 1412.835000 0.630000 ;
      RECT 1406.275000 0.000000 1409.345000 0.630000 ;
      RECT 1402.790000 0.000000 1405.855000 0.630000 ;
      RECT 1399.300000 0.000000 1402.370000 0.630000 ;
      RECT 1395.810000 0.000000 1398.880000 0.630000 ;
      RECT 1392.320000 0.000000 1395.390000 0.630000 ;
      RECT 1388.830000 0.000000 1391.900000 0.630000 ;
      RECT 1385.345000 0.000000 1388.410000 0.630000 ;
      RECT 1381.855000 0.000000 1384.925000 0.630000 ;
      RECT 1378.365000 0.000000 1381.435000 0.630000 ;
      RECT 1374.875000 0.000000 1377.945000 0.630000 ;
      RECT 1371.385000 0.000000 1374.455000 0.630000 ;
      RECT 1367.900000 0.000000 1370.965000 0.630000 ;
      RECT 1364.410000 0.000000 1367.480000 0.630000 ;
      RECT 1360.920000 0.000000 1363.990000 0.630000 ;
      RECT 1357.430000 0.000000 1360.500000 0.630000 ;
      RECT 1353.940000 0.000000 1357.010000 0.630000 ;
      RECT 1350.455000 0.000000 1353.520000 0.630000 ;
      RECT 1346.965000 0.000000 1350.035000 0.630000 ;
      RECT 1343.475000 0.000000 1346.545000 0.630000 ;
      RECT 1339.985000 0.000000 1343.055000 0.630000 ;
      RECT 1336.495000 0.000000 1339.565000 0.630000 ;
      RECT 1333.010000 0.000000 1336.075000 0.630000 ;
      RECT 1329.520000 0.000000 1332.590000 0.630000 ;
      RECT 1326.030000 0.000000 1329.100000 0.630000 ;
      RECT 1322.540000 0.000000 1325.610000 0.630000 ;
      RECT 1319.050000 0.000000 1322.120000 0.630000 ;
      RECT 1315.565000 0.000000 1318.630000 0.630000 ;
      RECT 1312.075000 0.000000 1315.145000 0.630000 ;
      RECT 1308.585000 0.000000 1311.655000 0.630000 ;
      RECT 1305.095000 0.000000 1308.165000 0.630000 ;
      RECT 1301.605000 0.000000 1304.675000 0.630000 ;
      RECT 1298.120000 0.000000 1301.185000 0.630000 ;
      RECT 1294.630000 0.000000 1297.700000 0.630000 ;
      RECT 1291.140000 0.000000 1294.210000 0.630000 ;
      RECT 1287.650000 0.000000 1290.720000 0.630000 ;
      RECT 1284.160000 0.000000 1287.230000 0.630000 ;
      RECT 1280.675000 0.000000 1283.740000 0.630000 ;
      RECT 1277.185000 0.000000 1280.255000 0.630000 ;
      RECT 1273.695000 0.000000 1276.765000 0.630000 ;
      RECT 1270.205000 0.000000 1273.275000 0.630000 ;
      RECT 1266.715000 0.000000 1269.785000 0.630000 ;
      RECT 1263.230000 0.000000 1266.295000 0.630000 ;
      RECT 1259.740000 0.000000 1262.810000 0.630000 ;
      RECT 1256.250000 0.000000 1259.320000 0.630000 ;
      RECT 1252.760000 0.000000 1255.830000 0.630000 ;
      RECT 1249.270000 0.000000 1252.340000 0.630000 ;
      RECT 1245.785000 0.000000 1248.850000 0.630000 ;
      RECT 1242.295000 0.000000 1245.365000 0.630000 ;
      RECT 1238.805000 0.000000 1241.875000 0.630000 ;
      RECT 1235.315000 0.000000 1238.385000 0.630000 ;
      RECT 1231.825000 0.000000 1234.895000 0.630000 ;
      RECT 1228.340000 0.000000 1231.405000 0.630000 ;
      RECT 1224.850000 0.000000 1227.920000 0.630000 ;
      RECT 1221.360000 0.000000 1224.430000 0.630000 ;
      RECT 1217.870000 0.000000 1220.940000 0.630000 ;
      RECT 1214.380000 0.000000 1217.450000 0.630000 ;
      RECT 1210.895000 0.000000 1213.960000 0.630000 ;
      RECT 1207.405000 0.000000 1210.475000 0.630000 ;
      RECT 1203.915000 0.000000 1206.985000 0.630000 ;
      RECT 1200.425000 0.000000 1203.495000 0.630000 ;
      RECT 1196.935000 0.000000 1200.005000 0.630000 ;
      RECT 1193.450000 0.000000 1196.515000 0.630000 ;
      RECT 1189.960000 0.000000 1193.030000 0.630000 ;
      RECT 1186.470000 0.000000 1189.540000 0.630000 ;
      RECT 1182.980000 0.000000 1186.050000 0.630000 ;
      RECT 1179.490000 0.000000 1182.560000 0.630000 ;
      RECT 1176.005000 0.000000 1179.070000 0.630000 ;
      RECT 1172.515000 0.000000 1175.585000 0.630000 ;
      RECT 1169.025000 0.000000 1172.095000 0.630000 ;
      RECT 1165.535000 0.000000 1168.605000 0.630000 ;
      RECT 1162.045000 0.000000 1165.115000 0.630000 ;
      RECT 1158.560000 0.000000 1161.625000 0.630000 ;
      RECT 1155.070000 0.000000 1158.140000 0.630000 ;
      RECT 1151.580000 0.000000 1154.650000 0.630000 ;
      RECT 1148.090000 0.000000 1151.160000 0.630000 ;
      RECT 1144.600000 0.000000 1147.670000 0.630000 ;
      RECT 1141.115000 0.000000 1144.180000 0.630000 ;
      RECT 1137.625000 0.000000 1140.695000 0.630000 ;
      RECT 1134.135000 0.000000 1137.205000 0.630000 ;
      RECT 1130.645000 0.000000 1133.715000 0.630000 ;
      RECT 1127.155000 0.000000 1130.225000 0.630000 ;
      RECT 1123.670000 0.000000 1126.735000 0.630000 ;
      RECT 1120.180000 0.000000 1123.250000 0.630000 ;
      RECT 1116.690000 0.000000 1119.760000 0.630000 ;
      RECT 1113.200000 0.000000 1116.270000 0.630000 ;
      RECT 1109.710000 0.000000 1112.780000 0.630000 ;
      RECT 1106.225000 0.000000 1109.290000 0.630000 ;
      RECT 1102.735000 0.000000 1105.805000 0.630000 ;
      RECT 1099.245000 0.000000 1102.315000 0.630000 ;
      RECT 1095.755000 0.000000 1098.825000 0.630000 ;
      RECT 1092.265000 0.000000 1095.335000 0.630000 ;
      RECT 1088.780000 0.000000 1091.845000 0.630000 ;
      RECT 1085.290000 0.000000 1088.360000 0.630000 ;
      RECT 1081.800000 0.000000 1084.870000 0.630000 ;
      RECT 1078.310000 0.000000 1081.380000 0.630000 ;
      RECT 1074.820000 0.000000 1077.890000 0.630000 ;
      RECT 1071.335000 0.000000 1074.400000 0.630000 ;
      RECT 1067.845000 0.000000 1070.915000 0.630000 ;
      RECT 1064.355000 0.000000 1067.425000 0.630000 ;
      RECT 1060.865000 0.000000 1063.935000 0.630000 ;
      RECT 1057.375000 0.000000 1060.445000 0.630000 ;
      RECT 1053.890000 0.000000 1056.955000 0.630000 ;
      RECT 1050.400000 0.000000 1053.470000 0.630000 ;
      RECT 1046.910000 0.000000 1049.980000 0.630000 ;
      RECT 1043.420000 0.000000 1046.490000 0.630000 ;
      RECT 1039.930000 0.000000 1043.000000 0.630000 ;
      RECT 1036.445000 0.000000 1039.510000 0.630000 ;
      RECT 1032.955000 0.000000 1036.025000 0.630000 ;
      RECT 1029.465000 0.000000 1032.535000 0.630000 ;
      RECT 1025.975000 0.000000 1029.045000 0.630000 ;
      RECT 1022.485000 0.000000 1025.555000 0.630000 ;
      RECT 1019.000000 0.000000 1022.065000 0.630000 ;
      RECT 1015.510000 0.000000 1018.580000 0.630000 ;
      RECT 1012.020000 0.000000 1015.090000 0.630000 ;
      RECT 1008.530000 0.000000 1011.600000 0.630000 ;
      RECT 1005.040000 0.000000 1008.110000 0.630000 ;
      RECT 1001.555000 0.000000 1004.620000 0.630000 ;
      RECT 998.065000 0.000000 1001.135000 0.630000 ;
      RECT 994.575000 0.000000 997.645000 0.630000 ;
      RECT 991.085000 0.000000 994.155000 0.630000 ;
      RECT 987.595000 0.000000 990.665000 0.630000 ;
      RECT 984.110000 0.000000 987.175000 0.630000 ;
      RECT 980.620000 0.000000 983.690000 0.630000 ;
      RECT 977.130000 0.000000 980.200000 0.630000 ;
      RECT 973.640000 0.000000 976.710000 0.630000 ;
      RECT 970.150000 0.000000 973.220000 0.630000 ;
      RECT 966.665000 0.000000 969.730000 0.630000 ;
      RECT 963.175000 0.000000 966.245000 0.630000 ;
      RECT 959.685000 0.000000 962.755000 0.630000 ;
      RECT 956.195000 0.000000 959.265000 0.630000 ;
      RECT 952.705000 0.000000 955.775000 0.630000 ;
      RECT 949.220000 0.000000 952.285000 0.630000 ;
      RECT 945.730000 0.000000 948.800000 0.630000 ;
      RECT 942.240000 0.000000 945.310000 0.630000 ;
      RECT 938.750000 0.000000 941.820000 0.630000 ;
      RECT 935.260000 0.000000 938.330000 0.630000 ;
      RECT 931.775000 0.000000 934.840000 0.630000 ;
      RECT 928.285000 0.000000 931.355000 0.630000 ;
      RECT 924.795000 0.000000 927.865000 0.630000 ;
      RECT 921.305000 0.000000 924.375000 0.630000 ;
      RECT 917.815000 0.000000 920.885000 0.630000 ;
      RECT 914.330000 0.000000 917.395000 0.630000 ;
      RECT 910.840000 0.000000 913.910000 0.630000 ;
      RECT 907.350000 0.000000 910.420000 0.630000 ;
      RECT 903.860000 0.000000 906.930000 0.630000 ;
      RECT 900.370000 0.000000 903.440000 0.630000 ;
      RECT 896.885000 0.000000 899.950000 0.630000 ;
      RECT 893.395000 0.000000 896.465000 0.630000 ;
      RECT 889.905000 0.000000 892.975000 0.630000 ;
      RECT 886.415000 0.000000 889.485000 0.630000 ;
      RECT 882.925000 0.000000 885.995000 0.630000 ;
      RECT 879.440000 0.000000 882.505000 0.630000 ;
      RECT 875.950000 0.000000 879.020000 0.630000 ;
      RECT 872.460000 0.000000 875.530000 0.630000 ;
      RECT 868.970000 0.000000 872.040000 0.630000 ;
      RECT 865.480000 0.000000 868.550000 0.630000 ;
      RECT 861.995000 0.000000 865.060000 0.630000 ;
      RECT 858.505000 0.000000 861.575000 0.630000 ;
      RECT 855.015000 0.000000 858.085000 0.630000 ;
      RECT 851.525000 0.000000 854.595000 0.630000 ;
      RECT 848.035000 0.000000 851.105000 0.630000 ;
      RECT 844.550000 0.000000 847.615000 0.630000 ;
      RECT 841.060000 0.000000 844.130000 0.630000 ;
      RECT 837.570000 0.000000 840.640000 0.630000 ;
      RECT 834.080000 0.000000 837.150000 0.630000 ;
      RECT 830.590000 0.000000 833.660000 0.630000 ;
      RECT 827.105000 0.000000 830.170000 0.630000 ;
      RECT 823.615000 0.000000 826.685000 0.630000 ;
      RECT 820.125000 0.000000 823.195000 0.630000 ;
      RECT 816.635000 0.000000 819.705000 0.630000 ;
      RECT 813.145000 0.000000 816.215000 0.630000 ;
      RECT 809.660000 0.000000 812.725000 0.630000 ;
      RECT 806.170000 0.000000 809.240000 0.630000 ;
      RECT 802.680000 0.000000 805.750000 0.630000 ;
      RECT 799.190000 0.000000 802.260000 0.630000 ;
      RECT 795.700000 0.000000 798.770000 0.630000 ;
      RECT 792.215000 0.000000 795.280000 0.630000 ;
      RECT 788.725000 0.000000 791.795000 0.630000 ;
      RECT 785.235000 0.000000 788.305000 0.630000 ;
      RECT 781.745000 0.000000 784.815000 0.630000 ;
      RECT 778.255000 0.000000 781.325000 0.630000 ;
      RECT 774.770000 0.000000 777.835000 0.630000 ;
      RECT 771.280000 0.000000 774.350000 0.630000 ;
      RECT 767.790000 0.000000 770.860000 0.630000 ;
      RECT 764.300000 0.000000 767.370000 0.630000 ;
      RECT 760.810000 0.000000 763.880000 0.630000 ;
      RECT 757.325000 0.000000 760.390000 0.630000 ;
      RECT 753.835000 0.000000 756.905000 0.630000 ;
      RECT 750.345000 0.000000 753.415000 0.630000 ;
      RECT 746.855000 0.000000 749.925000 0.630000 ;
      RECT 743.365000 0.000000 746.435000 0.630000 ;
      RECT 739.880000 0.000000 742.945000 0.630000 ;
      RECT 736.390000 0.000000 739.460000 0.630000 ;
      RECT 732.900000 0.000000 735.970000 0.630000 ;
      RECT 729.410000 0.000000 732.480000 0.630000 ;
      RECT 725.920000 0.000000 728.990000 0.630000 ;
      RECT 722.435000 0.000000 725.500000 0.630000 ;
      RECT 718.945000 0.000000 722.015000 0.630000 ;
      RECT 715.455000 0.000000 718.525000 0.630000 ;
      RECT 711.965000 0.000000 715.035000 0.630000 ;
      RECT 708.475000 0.000000 711.545000 0.630000 ;
      RECT 704.990000 0.000000 708.055000 0.630000 ;
      RECT 701.500000 0.000000 704.570000 0.630000 ;
      RECT 698.010000 0.000000 701.080000 0.630000 ;
      RECT 694.520000 0.000000 697.590000 0.630000 ;
      RECT 691.030000 0.000000 694.100000 0.630000 ;
      RECT 687.545000 0.000000 690.610000 0.630000 ;
      RECT 684.055000 0.000000 687.125000 0.630000 ;
      RECT 680.565000 0.000000 683.635000 0.630000 ;
      RECT 677.075000 0.000000 680.145000 0.630000 ;
      RECT 673.585000 0.000000 676.655000 0.630000 ;
      RECT 670.100000 0.000000 673.165000 0.630000 ;
      RECT 666.610000 0.000000 669.680000 0.630000 ;
      RECT 663.120000 0.000000 666.190000 0.630000 ;
      RECT 659.630000 0.000000 662.700000 0.630000 ;
      RECT 656.140000 0.000000 659.210000 0.630000 ;
      RECT 652.655000 0.000000 655.720000 0.630000 ;
      RECT 649.165000 0.000000 652.235000 0.630000 ;
      RECT 645.675000 0.000000 648.745000 0.630000 ;
      RECT 642.185000 0.000000 645.255000 0.630000 ;
      RECT 638.695000 0.000000 641.765000 0.630000 ;
      RECT 635.210000 0.000000 638.275000 0.630000 ;
      RECT 631.720000 0.000000 634.790000 0.630000 ;
      RECT 628.230000 0.000000 631.300000 0.630000 ;
      RECT 624.740000 0.000000 627.810000 0.630000 ;
      RECT 621.250000 0.000000 624.320000 0.630000 ;
      RECT 617.765000 0.000000 620.830000 0.630000 ;
      RECT 614.275000 0.000000 617.345000 0.630000 ;
      RECT 610.785000 0.000000 613.855000 0.630000 ;
      RECT 607.295000 0.000000 610.365000 0.630000 ;
      RECT 603.805000 0.000000 606.875000 0.630000 ;
      RECT 600.320000 0.000000 603.385000 0.630000 ;
      RECT 596.830000 0.000000 599.900000 0.630000 ;
      RECT 593.340000 0.000000 596.410000 0.630000 ;
      RECT 589.850000 0.000000 592.920000 0.630000 ;
      RECT 586.360000 0.000000 589.430000 0.630000 ;
      RECT 582.875000 0.000000 585.940000 0.630000 ;
      RECT 579.385000 0.000000 582.455000 0.630000 ;
      RECT 575.895000 0.000000 578.965000 0.630000 ;
      RECT 572.405000 0.000000 575.475000 0.630000 ;
      RECT 568.915000 0.000000 571.985000 0.630000 ;
      RECT 565.430000 0.000000 568.495000 0.630000 ;
      RECT 561.940000 0.000000 565.010000 0.630000 ;
      RECT 558.450000 0.000000 561.520000 0.630000 ;
      RECT 554.960000 0.000000 558.030000 0.630000 ;
      RECT 551.470000 0.000000 554.540000 0.630000 ;
      RECT 547.985000 0.000000 551.050000 0.630000 ;
      RECT 544.495000 0.000000 547.565000 0.630000 ;
      RECT 541.005000 0.000000 544.075000 0.630000 ;
      RECT 537.515000 0.000000 540.585000 0.630000 ;
      RECT 534.025000 0.000000 537.095000 0.630000 ;
      RECT 530.540000 0.000000 533.605000 0.630000 ;
      RECT 527.050000 0.000000 530.120000 0.630000 ;
      RECT 523.560000 0.000000 526.630000 0.630000 ;
      RECT 520.070000 0.000000 523.140000 0.630000 ;
      RECT 516.580000 0.000000 519.650000 0.630000 ;
      RECT 513.095000 0.000000 516.160000 0.630000 ;
      RECT 509.605000 0.000000 512.675000 0.630000 ;
      RECT 506.115000 0.000000 509.185000 0.630000 ;
      RECT 502.625000 0.000000 505.695000 0.630000 ;
      RECT 499.135000 0.000000 502.205000 0.630000 ;
      RECT 495.650000 0.000000 498.715000 0.630000 ;
      RECT 492.160000 0.000000 495.230000 0.630000 ;
      RECT 488.670000 0.000000 491.740000 0.630000 ;
      RECT 485.180000 0.000000 488.250000 0.630000 ;
      RECT 481.690000 0.000000 484.760000 0.630000 ;
      RECT 478.205000 0.000000 481.270000 0.630000 ;
      RECT 474.715000 0.000000 477.785000 0.630000 ;
      RECT 471.225000 0.000000 474.295000 0.630000 ;
      RECT 467.735000 0.000000 470.805000 0.630000 ;
      RECT 464.245000 0.000000 467.315000 0.630000 ;
      RECT 460.760000 0.000000 463.825000 0.630000 ;
      RECT 457.270000 0.000000 460.340000 0.630000 ;
      RECT 453.780000 0.000000 456.850000 0.630000 ;
      RECT 450.290000 0.000000 453.360000 0.630000 ;
      RECT 446.800000 0.000000 449.870000 0.630000 ;
      RECT 443.315000 0.000000 446.380000 0.630000 ;
      RECT 439.825000 0.000000 442.895000 0.630000 ;
      RECT 436.335000 0.000000 439.405000 0.630000 ;
      RECT 432.845000 0.000000 435.915000 0.630000 ;
      RECT 429.355000 0.000000 432.425000 0.630000 ;
      RECT 425.870000 0.000000 428.935000 0.630000 ;
      RECT 422.380000 0.000000 425.450000 0.630000 ;
      RECT 418.890000 0.000000 421.960000 0.630000 ;
      RECT 415.400000 0.000000 418.470000 0.630000 ;
      RECT 411.910000 0.000000 414.980000 0.630000 ;
      RECT 408.425000 0.000000 411.490000 0.630000 ;
      RECT 404.935000 0.000000 408.005000 0.630000 ;
      RECT 401.445000 0.000000 404.515000 0.630000 ;
      RECT 397.955000 0.000000 401.025000 0.630000 ;
      RECT 394.465000 0.000000 397.535000 0.630000 ;
      RECT 390.980000 0.000000 394.045000 0.630000 ;
      RECT 387.490000 0.000000 390.560000 0.630000 ;
      RECT 384.000000 0.000000 387.070000 0.630000 ;
      RECT 380.510000 0.000000 383.580000 0.630000 ;
      RECT 377.020000 0.000000 380.090000 0.630000 ;
      RECT 373.535000 0.000000 376.600000 0.630000 ;
      RECT 370.045000 0.000000 373.115000 0.630000 ;
      RECT 366.555000 0.000000 369.625000 0.630000 ;
      RECT 363.065000 0.000000 366.135000 0.630000 ;
      RECT 359.575000 0.000000 362.645000 0.630000 ;
      RECT 356.090000 0.000000 359.155000 0.630000 ;
      RECT 352.600000 0.000000 355.670000 0.630000 ;
      RECT 349.110000 0.000000 352.180000 0.630000 ;
      RECT 345.620000 0.000000 348.690000 0.630000 ;
      RECT 342.130000 0.000000 345.200000 0.630000 ;
      RECT 338.645000 0.000000 341.710000 0.630000 ;
      RECT 335.155000 0.000000 338.225000 0.630000 ;
      RECT 331.665000 0.000000 334.735000 0.630000 ;
      RECT 328.175000 0.000000 331.245000 0.630000 ;
      RECT 324.685000 0.000000 327.755000 0.630000 ;
      RECT 321.200000 0.000000 324.265000 0.630000 ;
      RECT 317.710000 0.000000 320.780000 0.630000 ;
      RECT 314.220000 0.000000 317.290000 0.630000 ;
      RECT 310.730000 0.000000 313.800000 0.630000 ;
      RECT 307.240000 0.000000 310.310000 0.630000 ;
      RECT 303.755000 0.000000 306.820000 0.630000 ;
      RECT 300.265000 0.000000 303.335000 0.630000 ;
      RECT 296.775000 0.000000 299.845000 0.630000 ;
      RECT 293.285000 0.000000 296.355000 0.630000 ;
      RECT 289.795000 0.000000 292.865000 0.630000 ;
      RECT 286.310000 0.000000 289.375000 0.630000 ;
      RECT 282.820000 0.000000 285.890000 0.630000 ;
      RECT 279.330000 0.000000 282.400000 0.630000 ;
      RECT 275.840000 0.000000 278.910000 0.630000 ;
      RECT 272.350000 0.000000 275.420000 0.630000 ;
      RECT 268.865000 0.000000 271.930000 0.630000 ;
      RECT 265.375000 0.000000 268.445000 0.630000 ;
      RECT 261.885000 0.000000 264.955000 0.630000 ;
      RECT 258.395000 0.000000 261.465000 0.630000 ;
      RECT 254.905000 0.000000 257.975000 0.630000 ;
      RECT 251.420000 0.000000 254.485000 0.630000 ;
      RECT 247.930000 0.000000 251.000000 0.630000 ;
      RECT 244.440000 0.000000 247.510000 0.630000 ;
      RECT 240.950000 0.000000 244.020000 0.630000 ;
      RECT 237.460000 0.000000 240.530000 0.630000 ;
      RECT 233.975000 0.000000 237.040000 0.630000 ;
      RECT 230.485000 0.000000 233.555000 0.630000 ;
      RECT 226.995000 0.000000 230.065000 0.630000 ;
      RECT 223.505000 0.000000 226.575000 0.630000 ;
      RECT 220.015000 0.000000 223.085000 0.630000 ;
      RECT 216.530000 0.000000 219.595000 0.630000 ;
      RECT 213.040000 0.000000 216.110000 0.630000 ;
      RECT 209.550000 0.000000 212.620000 0.630000 ;
      RECT 206.060000 0.000000 209.130000 0.630000 ;
      RECT 202.570000 0.000000 205.640000 0.630000 ;
      RECT 199.085000 0.000000 202.150000 0.630000 ;
      RECT 195.595000 0.000000 198.665000 0.630000 ;
      RECT 192.105000 0.000000 195.175000 0.630000 ;
      RECT 188.615000 0.000000 191.685000 0.630000 ;
      RECT 185.125000 0.000000 188.195000 0.630000 ;
      RECT 181.640000 0.000000 184.705000 0.630000 ;
      RECT 178.150000 0.000000 181.220000 0.630000 ;
      RECT 174.660000 0.000000 177.730000 0.630000 ;
      RECT 171.170000 0.000000 174.240000 0.630000 ;
      RECT 167.680000 0.000000 170.750000 0.630000 ;
      RECT 164.195000 0.000000 167.260000 0.630000 ;
      RECT 160.705000 0.000000 163.775000 0.630000 ;
      RECT 157.215000 0.000000 160.285000 0.630000 ;
      RECT 153.725000 0.000000 156.795000 0.630000 ;
      RECT 150.235000 0.000000 153.305000 0.630000 ;
      RECT 146.750000 0.000000 149.815000 0.630000 ;
      RECT 143.260000 0.000000 146.330000 0.630000 ;
      RECT 139.770000 0.000000 142.840000 0.630000 ;
      RECT 136.280000 0.000000 139.350000 0.630000 ;
      RECT 132.790000 0.000000 135.860000 0.630000 ;
      RECT 129.305000 0.000000 132.370000 0.630000 ;
      RECT 125.815000 0.000000 128.885000 0.630000 ;
      RECT 122.325000 0.000000 125.395000 0.630000 ;
      RECT 118.835000 0.000000 121.905000 0.630000 ;
      RECT 115.345000 0.000000 118.415000 0.630000 ;
      RECT 111.860000 0.000000 114.925000 0.630000 ;
      RECT 108.370000 0.000000 111.440000 0.630000 ;
      RECT 104.880000 0.000000 107.950000 0.630000 ;
      RECT 101.390000 0.000000 104.460000 0.630000 ;
      RECT 97.900000 0.000000 100.970000 0.630000 ;
      RECT 94.415000 0.000000 97.480000 0.630000 ;
      RECT 90.925000 0.000000 93.995000 0.630000 ;
      RECT 87.435000 0.000000 90.505000 0.630000 ;
      RECT 83.945000 0.000000 87.015000 0.630000 ;
      RECT 80.455000 0.000000 83.525000 0.630000 ;
      RECT 76.970000 0.000000 80.035000 0.630000 ;
      RECT 73.480000 0.000000 76.550000 0.630000 ;
      RECT 69.990000 0.000000 73.060000 0.630000 ;
      RECT 66.500000 0.000000 69.570000 0.630000 ;
      RECT 63.010000 0.000000 66.080000 0.630000 ;
      RECT 59.525000 0.000000 62.590000 0.630000 ;
      RECT 56.035000 0.000000 59.105000 0.630000 ;
      RECT 52.545000 0.000000 55.615000 0.630000 ;
      RECT 49.055000 0.000000 52.125000 0.630000 ;
      RECT 45.565000 0.000000 48.635000 0.630000 ;
      RECT 42.080000 0.000000 45.145000 0.630000 ;
      RECT 38.590000 0.000000 41.660000 0.630000 ;
      RECT 35.100000 0.000000 38.170000 0.630000 ;
      RECT 31.610000 0.000000 34.680000 0.630000 ;
      RECT 28.120000 0.000000 31.190000 0.630000 ;
      RECT 24.635000 0.000000 27.700000 0.630000 ;
      RECT 21.145000 0.000000 24.215000 0.630000 ;
      RECT 17.655000 0.000000 20.725000 0.630000 ;
      RECT 14.165000 0.000000 17.235000 0.630000 ;
      RECT 10.675000 0.000000 13.745000 0.630000 ;
      RECT 7.190000 0.000000 10.255000 0.630000 ;
      RECT 3.700000 0.000000 6.770000 0.630000 ;
      RECT 1.820000 0.000000 3.280000 0.630000 ;
      RECT 0.000000 0.000000 1.400000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 1465.940000 1720.400000 1469.820000 ;
      RECT 1.100000 1465.330000 1720.400000 1465.940000 ;
      RECT 1.100000 1465.040000 1719.300000 1465.330000 ;
      RECT 0.000000 1464.430000 1719.300000 1465.040000 ;
      RECT 0.000000 1442.515000 1720.400000 1464.430000 ;
      RECT 1.100000 1441.965000 1720.400000 1442.515000 ;
      RECT 1.100000 1441.615000 1719.300000 1441.965000 ;
      RECT 0.000000 1441.065000 1719.300000 1441.615000 ;
      RECT 0.000000 1414.780000 1720.400000 1441.065000 ;
      RECT 1.100000 1413.880000 1720.400000 1414.780000 ;
      RECT 0.000000 1413.700000 1720.400000 1413.880000 ;
      RECT 0.000000 1412.800000 1719.300000 1413.700000 ;
      RECT 0.000000 1387.050000 1720.400000 1412.800000 ;
      RECT 1.100000 1386.150000 1720.400000 1387.050000 ;
      RECT 0.000000 1385.435000 1720.400000 1386.150000 ;
      RECT 0.000000 1384.535000 1719.300000 1385.435000 ;
      RECT 0.000000 1359.320000 1720.400000 1384.535000 ;
      RECT 1.100000 1358.420000 1720.400000 1359.320000 ;
      RECT 0.000000 1357.170000 1720.400000 1358.420000 ;
      RECT 0.000000 1356.270000 1719.300000 1357.170000 ;
      RECT 0.000000 1331.585000 1720.400000 1356.270000 ;
      RECT 1.100000 1330.685000 1720.400000 1331.585000 ;
      RECT 0.000000 1328.905000 1720.400000 1330.685000 ;
      RECT 0.000000 1328.005000 1719.300000 1328.905000 ;
      RECT 0.000000 1303.855000 1720.400000 1328.005000 ;
      RECT 1.100000 1302.955000 1720.400000 1303.855000 ;
      RECT 0.000000 1300.640000 1720.400000 1302.955000 ;
      RECT 0.000000 1299.740000 1719.300000 1300.640000 ;
      RECT 0.000000 1276.120000 1720.400000 1299.740000 ;
      RECT 1.100000 1275.220000 1720.400000 1276.120000 ;
      RECT 0.000000 1272.375000 1720.400000 1275.220000 ;
      RECT 0.000000 1271.475000 1719.300000 1272.375000 ;
      RECT 0.000000 1248.390000 1720.400000 1271.475000 ;
      RECT 1.100000 1247.490000 1720.400000 1248.390000 ;
      RECT 0.000000 1244.110000 1720.400000 1247.490000 ;
      RECT 0.000000 1243.210000 1719.300000 1244.110000 ;
      RECT 0.000000 1220.660000 1720.400000 1243.210000 ;
      RECT 1.100000 1219.760000 1720.400000 1220.660000 ;
      RECT 0.000000 1215.845000 1720.400000 1219.760000 ;
      RECT 0.000000 1214.945000 1719.300000 1215.845000 ;
      RECT 0.000000 1192.925000 1720.400000 1214.945000 ;
      RECT 1.100000 1192.025000 1720.400000 1192.925000 ;
      RECT 0.000000 1187.580000 1720.400000 1192.025000 ;
      RECT 0.000000 1186.680000 1719.300000 1187.580000 ;
      RECT 0.000000 1165.195000 1720.400000 1186.680000 ;
      RECT 1.100000 1164.295000 1720.400000 1165.195000 ;
      RECT 0.000000 1159.315000 1720.400000 1164.295000 ;
      RECT 0.000000 1158.415000 1719.300000 1159.315000 ;
      RECT 0.000000 1137.460000 1720.400000 1158.415000 ;
      RECT 1.100000 1136.560000 1720.400000 1137.460000 ;
      RECT 0.000000 1131.050000 1720.400000 1136.560000 ;
      RECT 0.000000 1130.150000 1719.300000 1131.050000 ;
      RECT 0.000000 1109.730000 1720.400000 1130.150000 ;
      RECT 1.100000 1108.830000 1720.400000 1109.730000 ;
      RECT 0.000000 1102.785000 1720.400000 1108.830000 ;
      RECT 0.000000 1101.885000 1719.300000 1102.785000 ;
      RECT 0.000000 1082.000000 1720.400000 1101.885000 ;
      RECT 1.100000 1081.100000 1720.400000 1082.000000 ;
      RECT 0.000000 1074.520000 1720.400000 1081.100000 ;
      RECT 0.000000 1073.620000 1719.300000 1074.520000 ;
      RECT 0.000000 1054.265000 1720.400000 1073.620000 ;
      RECT 1.100000 1053.365000 1720.400000 1054.265000 ;
      RECT 0.000000 1046.255000 1720.400000 1053.365000 ;
      RECT 0.000000 1045.355000 1719.300000 1046.255000 ;
      RECT 0.000000 1026.535000 1720.400000 1045.355000 ;
      RECT 1.100000 1025.635000 1720.400000 1026.535000 ;
      RECT 0.000000 1017.990000 1720.400000 1025.635000 ;
      RECT 0.000000 1017.090000 1719.300000 1017.990000 ;
      RECT 0.000000 998.800000 1720.400000 1017.090000 ;
      RECT 1.100000 997.900000 1720.400000 998.800000 ;
      RECT 0.000000 989.725000 1720.400000 997.900000 ;
      RECT 0.000000 988.825000 1719.300000 989.725000 ;
      RECT 0.000000 971.070000 1720.400000 988.825000 ;
      RECT 1.100000 970.170000 1720.400000 971.070000 ;
      RECT 0.000000 961.460000 1720.400000 970.170000 ;
      RECT 0.000000 960.560000 1719.300000 961.460000 ;
      RECT 0.000000 943.340000 1720.400000 960.560000 ;
      RECT 1.100000 942.440000 1720.400000 943.340000 ;
      RECT 0.000000 933.195000 1720.400000 942.440000 ;
      RECT 0.000000 932.295000 1719.300000 933.195000 ;
      RECT 0.000000 915.605000 1720.400000 932.295000 ;
      RECT 1.100000 914.705000 1720.400000 915.605000 ;
      RECT 0.000000 904.930000 1720.400000 914.705000 ;
      RECT 0.000000 904.030000 1719.300000 904.930000 ;
      RECT 0.000000 887.875000 1720.400000 904.030000 ;
      RECT 1.100000 886.975000 1720.400000 887.875000 ;
      RECT 0.000000 876.665000 1720.400000 886.975000 ;
      RECT 0.000000 875.765000 1719.300000 876.665000 ;
      RECT 0.000000 860.140000 1720.400000 875.765000 ;
      RECT 1.100000 859.240000 1720.400000 860.140000 ;
      RECT 0.000000 848.400000 1720.400000 859.240000 ;
      RECT 0.000000 847.500000 1719.300000 848.400000 ;
      RECT 0.000000 832.410000 1720.400000 847.500000 ;
      RECT 1.100000 831.510000 1720.400000 832.410000 ;
      RECT 0.000000 820.135000 1720.400000 831.510000 ;
      RECT 0.000000 819.235000 1719.300000 820.135000 ;
      RECT 0.000000 804.680000 1720.400000 819.235000 ;
      RECT 1.100000 803.780000 1720.400000 804.680000 ;
      RECT 0.000000 791.870000 1720.400000 803.780000 ;
      RECT 0.000000 790.970000 1719.300000 791.870000 ;
      RECT 0.000000 776.945000 1720.400000 790.970000 ;
      RECT 1.100000 776.045000 1720.400000 776.945000 ;
      RECT 0.000000 763.605000 1720.400000 776.045000 ;
      RECT 0.000000 762.705000 1719.300000 763.605000 ;
      RECT 0.000000 749.215000 1720.400000 762.705000 ;
      RECT 1.100000 748.315000 1720.400000 749.215000 ;
      RECT 0.000000 735.340000 1720.400000 748.315000 ;
      RECT 0.000000 734.440000 1719.300000 735.340000 ;
      RECT 0.000000 721.480000 1720.400000 734.440000 ;
      RECT 1.100000 720.580000 1720.400000 721.480000 ;
      RECT 0.000000 707.075000 1720.400000 720.580000 ;
      RECT 0.000000 706.175000 1719.300000 707.075000 ;
      RECT 0.000000 693.750000 1720.400000 706.175000 ;
      RECT 1.100000 692.850000 1720.400000 693.750000 ;
      RECT 0.000000 678.810000 1720.400000 692.850000 ;
      RECT 0.000000 677.910000 1719.300000 678.810000 ;
      RECT 0.000000 666.020000 1720.400000 677.910000 ;
      RECT 1.100000 665.120000 1720.400000 666.020000 ;
      RECT 0.000000 650.545000 1720.400000 665.120000 ;
      RECT 0.000000 649.645000 1719.300000 650.545000 ;
      RECT 0.000000 638.285000 1720.400000 649.645000 ;
      RECT 1.100000 637.385000 1720.400000 638.285000 ;
      RECT 0.000000 622.280000 1720.400000 637.385000 ;
      RECT 0.000000 621.380000 1719.300000 622.280000 ;
      RECT 0.000000 610.555000 1720.400000 621.380000 ;
      RECT 1.100000 609.655000 1720.400000 610.555000 ;
      RECT 0.000000 594.015000 1720.400000 609.655000 ;
      RECT 0.000000 593.115000 1719.300000 594.015000 ;
      RECT 0.000000 582.820000 1720.400000 593.115000 ;
      RECT 1.100000 581.920000 1720.400000 582.820000 ;
      RECT 0.000000 565.750000 1720.400000 581.920000 ;
      RECT 0.000000 564.850000 1719.300000 565.750000 ;
      RECT 0.000000 555.090000 1720.400000 564.850000 ;
      RECT 1.100000 554.190000 1720.400000 555.090000 ;
      RECT 0.000000 537.485000 1720.400000 554.190000 ;
      RECT 0.000000 536.585000 1719.300000 537.485000 ;
      RECT 0.000000 527.360000 1720.400000 536.585000 ;
      RECT 1.100000 526.460000 1720.400000 527.360000 ;
      RECT 0.000000 509.220000 1720.400000 526.460000 ;
      RECT 0.000000 508.320000 1719.300000 509.220000 ;
      RECT 0.000000 499.625000 1720.400000 508.320000 ;
      RECT 1.100000 498.725000 1720.400000 499.625000 ;
      RECT 0.000000 480.955000 1720.400000 498.725000 ;
      RECT 0.000000 480.055000 1719.300000 480.955000 ;
      RECT 0.000000 471.895000 1720.400000 480.055000 ;
      RECT 1.100000 470.995000 1720.400000 471.895000 ;
      RECT 0.000000 452.690000 1720.400000 470.995000 ;
      RECT 0.000000 451.790000 1719.300000 452.690000 ;
      RECT 0.000000 444.160000 1720.400000 451.790000 ;
      RECT 1.100000 443.260000 1720.400000 444.160000 ;
      RECT 0.000000 424.425000 1720.400000 443.260000 ;
      RECT 0.000000 423.525000 1719.300000 424.425000 ;
      RECT 0.000000 416.430000 1720.400000 423.525000 ;
      RECT 1.100000 415.530000 1720.400000 416.430000 ;
      RECT 0.000000 396.160000 1720.400000 415.530000 ;
      RECT 0.000000 395.260000 1719.300000 396.160000 ;
      RECT 0.000000 388.700000 1720.400000 395.260000 ;
      RECT 1.100000 387.800000 1720.400000 388.700000 ;
      RECT 0.000000 367.895000 1720.400000 387.800000 ;
      RECT 0.000000 366.995000 1719.300000 367.895000 ;
      RECT 0.000000 360.965000 1720.400000 366.995000 ;
      RECT 1.100000 360.065000 1720.400000 360.965000 ;
      RECT 0.000000 339.630000 1720.400000 360.065000 ;
      RECT 0.000000 338.730000 1719.300000 339.630000 ;
      RECT 0.000000 333.235000 1720.400000 338.730000 ;
      RECT 1.100000 332.335000 1720.400000 333.235000 ;
      RECT 0.000000 311.365000 1720.400000 332.335000 ;
      RECT 0.000000 310.465000 1719.300000 311.365000 ;
      RECT 0.000000 305.500000 1720.400000 310.465000 ;
      RECT 1.100000 304.600000 1720.400000 305.500000 ;
      RECT 0.000000 283.100000 1720.400000 304.600000 ;
      RECT 0.000000 282.200000 1719.300000 283.100000 ;
      RECT 0.000000 277.770000 1720.400000 282.200000 ;
      RECT 1.100000 276.870000 1720.400000 277.770000 ;
      RECT 0.000000 254.835000 1720.400000 276.870000 ;
      RECT 0.000000 253.935000 1719.300000 254.835000 ;
      RECT 0.000000 250.040000 1720.400000 253.935000 ;
      RECT 1.100000 249.140000 1720.400000 250.040000 ;
      RECT 0.000000 226.570000 1720.400000 249.140000 ;
      RECT 0.000000 225.670000 1719.300000 226.570000 ;
      RECT 0.000000 222.305000 1720.400000 225.670000 ;
      RECT 1.100000 221.405000 1720.400000 222.305000 ;
      RECT 0.000000 198.305000 1720.400000 221.405000 ;
      RECT 0.000000 197.405000 1719.300000 198.305000 ;
      RECT 0.000000 194.575000 1720.400000 197.405000 ;
      RECT 1.100000 193.675000 1720.400000 194.575000 ;
      RECT 0.000000 170.040000 1720.400000 193.675000 ;
      RECT 0.000000 169.140000 1719.300000 170.040000 ;
      RECT 0.000000 166.840000 1720.400000 169.140000 ;
      RECT 1.100000 165.940000 1720.400000 166.840000 ;
      RECT 0.000000 141.775000 1720.400000 165.940000 ;
      RECT 0.000000 140.875000 1719.300000 141.775000 ;
      RECT 0.000000 139.110000 1720.400000 140.875000 ;
      RECT 1.100000 138.210000 1720.400000 139.110000 ;
      RECT 0.000000 113.510000 1720.400000 138.210000 ;
      RECT 0.000000 112.610000 1719.300000 113.510000 ;
      RECT 0.000000 111.380000 1720.400000 112.610000 ;
      RECT 1.100000 110.480000 1720.400000 111.380000 ;
      RECT 0.000000 85.245000 1720.400000 110.480000 ;
      RECT 0.000000 84.345000 1719.300000 85.245000 ;
      RECT 0.000000 83.645000 1720.400000 84.345000 ;
      RECT 1.100000 82.745000 1720.400000 83.645000 ;
      RECT 0.000000 56.980000 1720.400000 82.745000 ;
      RECT 0.000000 56.080000 1719.300000 56.980000 ;
      RECT 0.000000 55.915000 1720.400000 56.080000 ;
      RECT 1.100000 55.015000 1720.400000 55.915000 ;
      RECT 0.000000 28.715000 1720.400000 55.015000 ;
      RECT 0.000000 28.180000 1719.300000 28.715000 ;
      RECT 1.100000 27.815000 1719.300000 28.180000 ;
      RECT 1.100000 27.280000 1720.400000 27.815000 ;
      RECT 0.000000 4.990000 1720.400000 27.280000 ;
      RECT 1.100000 4.380000 1720.400000 4.990000 ;
      RECT 1.100000 4.090000 1719.300000 4.380000 ;
      RECT 0.000000 3.480000 1719.300000 4.090000 ;
      RECT 0.000000 0.000000 1720.400000 3.480000 ;
    LAYER met4 ;
      RECT 0.000000 1468.020000 1720.400000 1469.820000 ;
      RECT 4.360000 1464.020000 1716.040000 1468.020000 ;
      RECT 1714.640000 5.630000 1716.040000 1464.020000 ;
      RECT 8.360000 5.630000 1712.040000 1464.020000 ;
      RECT 4.360000 5.630000 5.760000 1464.020000 ;
      RECT 1718.640000 1.630000 1720.400000 1468.020000 ;
      RECT 4.360000 1.630000 1716.040000 5.630000 ;
      RECT 0.000000 1.630000 1.760000 1468.020000 ;
      RECT 0.000000 0.000000 1720.400000 1.630000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
