##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Thu Dec 30 01:04:18 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 2220.420000 BY 2939.640000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.435000 0.000000 4.575000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.540000 0.000000 1.680000 0.490000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.240000 0.000000 468.380000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.535000 0.000000 157.675000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.745000 0.000000 472.885000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.740000 0.000000 463.880000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.235000 0.000000 459.375000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.735000 0.000000 454.875000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.230000 0.000000 450.370000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.630000 0.000000 301.770000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.130000 0.000000 297.270000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.625000 0.000000 292.765000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.120000 0.000000 288.260000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.620000 0.000000 283.760000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.115000 0.000000 279.255000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.615000 0.000000 274.755000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110000 0.000000 270.250000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.605000 0.000000 265.745000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.105000 0.000000 261.245000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.600000 0.000000 256.740000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.100000 0.000000 252.240000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.595000 0.000000 247.735000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.090000 0.000000 243.230000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.590000 0.000000 238.730000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.085000 0.000000 234.225000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.585000 0.000000 229.725000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.080000 0.000000 225.220000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.575000 0.000000 220.715000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.075000 0.000000 216.215000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.570000 0.000000 211.710000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.070000 0.000000 207.210000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.565000 0.000000 202.705000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.060000 0.000000 198.200000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.560000 0.000000 193.700000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.055000 0.000000 189.195000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.555000 0.000000 184.695000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.050000 0.000000 180.190000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.545000 0.000000 175.685000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.045000 0.000000 171.185000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.540000 0.000000 166.680000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.040000 0.000000 162.180000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.030000 0.000000 153.170000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.530000 0.000000 148.670000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.025000 0.000000 144.165000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.525000 0.000000 139.665000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.020000 0.000000 135.160000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.515000 0.000000 130.655000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.015000 0.000000 126.155000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.510000 0.000000 121.650000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.010000 0.000000 117.150000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.505000 0.000000 112.645000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.000000 0.000000 108.140000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.500000 0.000000 103.640000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.995000 0.000000 99.135000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.495000 0.000000 94.635000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.990000 0.000000 90.130000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.485000 0.000000 85.625000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.985000 0.000000 81.125000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.480000 0.000000 76.620000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.980000 0.000000 72.120000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.475000 0.000000 67.615000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.970000 0.000000 63.110000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.470000 0.000000 58.610000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.965000 0.000000 54.105000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.465000 0.000000 49.605000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.960000 0.000000 45.100000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.455000 0.000000 40.595000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.955000 0.000000 36.095000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.450000 0.000000 31.590000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.950000 0.000000 27.090000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.445000 0.000000 22.585000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.940000 0.000000 18.080000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.440000 0.000000 13.580000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.935000 0.000000 9.075000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.725000 0.000000 445.865000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.225000 0.000000 441.365000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.720000 0.000000 436.860000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.220000 0.000000 432.360000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.715000 0.000000 427.855000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.210000 0.000000 423.350000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.710000 0.000000 418.850000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.205000 0.000000 414.345000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.705000 0.000000 409.845000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.200000 0.000000 405.340000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.695000 0.000000 400.835000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.195000 0.000000 396.335000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.690000 0.000000 391.830000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.190000 0.000000 387.330000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.685000 0.000000 382.825000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.180000 0.000000 378.320000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.680000 0.000000 373.820000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.175000 0.000000 369.315000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.675000 0.000000 364.815000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.170000 0.000000 360.310000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.665000 0.000000 355.805000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.165000 0.000000 351.305000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.660000 0.000000 346.800000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.160000 0.000000 342.300000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.655000 0.000000 337.795000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.150000 0.000000 333.290000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.650000 0.000000 328.790000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.145000 0.000000 324.285000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.645000 0.000000 319.785000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.140000 0.000000 315.280000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.635000 0.000000 310.775000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.135000 0.000000 306.275000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.130000 0.000000 1049.270000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.625000 0.000000 1044.765000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.125000 0.000000 1040.265000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.620000 0.000000 1035.760000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.115000 0.000000 1031.255000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.615000 0.000000 1026.755000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.110000 0.000000 1022.250000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610000 0.000000 1017.750000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.105000 0.000000 1013.245000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.600000 0.000000 1008.740000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.100000 0.000000 1004.240000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.595000 0.000000 999.735000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.095000 0.000000 995.235000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.590000 0.000000 990.730000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.085000 0.000000 986.225000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.585000 0.000000 981.725000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.080000 0.000000 977.220000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.580000 0.000000 972.720000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.075000 0.000000 968.215000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.570000 0.000000 963.710000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.070000 0.000000 959.210000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.565000 0.000000 954.705000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.065000 0.000000 950.205000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.560000 0.000000 945.700000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.055000 0.000000 941.195000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.555000 0.000000 936.695000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050000 0.000000 932.190000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.550000 0.000000 927.690000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.045000 0.000000 923.185000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.540000 0.000000 918.680000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.040000 0.000000 914.180000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.535000 0.000000 909.675000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.035000 0.000000 905.175000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.530000 0.000000 900.670000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.025000 0.000000 896.165000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.525000 0.000000 891.665000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.020000 0.000000 887.160000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.520000 0.000000 882.660000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.015000 0.000000 878.155000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.510000 0.000000 873.650000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.010000 0.000000 869.150000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.505000 0.000000 864.645000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.005000 0.000000 860.145000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.500000 0.000000 855.640000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.995000 0.000000 851.135000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.495000 0.000000 846.635000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.990000 0.000000 842.130000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.490000 0.000000 837.630000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.985000 0.000000 833.125000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.480000 0.000000 828.620000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.980000 0.000000 824.120000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.475000 0.000000 819.615000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.975000 0.000000 815.115000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.470000 0.000000 810.610000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.965000 0.000000 806.105000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.465000 0.000000 801.605000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.960000 0.000000 797.100000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.460000 0.000000 792.600000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.955000 0.000000 788.095000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.450000 0.000000 783.590000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.950000 0.000000 779.090000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.445000 0.000000 774.585000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.945000 0.000000 770.085000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.440000 0.000000 765.580000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.935000 0.000000 761.075000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.435000 0.000000 756.575000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.930000 0.000000 752.070000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.430000 0.000000 747.570000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.925000 0.000000 743.065000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.420000 0.000000 738.560000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.920000 0.000000 734.060000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.415000 0.000000 729.555000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.915000 0.000000 725.055000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.410000 0.000000 720.550000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.905000 0.000000 716.045000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.405000 0.000000 711.545000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.900000 0.000000 707.040000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.400000 0.000000 702.540000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.895000 0.000000 698.035000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.390000 0.000000 693.530000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.890000 0.000000 689.030000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.385000 0.000000 684.525000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.885000 0.000000 680.025000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.380000 0.000000 675.520000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.875000 0.000000 671.015000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.375000 0.000000 666.515000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.870000 0.000000 662.010000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.370000 0.000000 657.510000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.865000 0.000000 653.005000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.360000 0.000000 648.500000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.860000 0.000000 644.000000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.355000 0.000000 639.495000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.855000 0.000000 634.995000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.350000 0.000000 630.490000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.845000 0.000000 625.985000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.345000 0.000000 621.485000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.840000 0.000000 616.980000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.340000 0.000000 612.480000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.835000 0.000000 607.975000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.330000 0.000000 603.470000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.830000 0.000000 598.970000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.325000 0.000000 594.465000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.825000 0.000000 589.965000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.320000 0.000000 585.460000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.815000 0.000000 580.955000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.315000 0.000000 576.455000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.810000 0.000000 571.950000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.310000 0.000000 567.450000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.805000 0.000000 562.945000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.300000 0.000000 558.440000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.800000 0.000000 553.940000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.295000 0.000000 549.435000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.795000 0.000000 544.935000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.290000 0.000000 540.430000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.785000 0.000000 535.925000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.285000 0.000000 531.425000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.780000 0.000000 526.920000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.280000 0.000000 522.420000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.775000 0.000000 517.915000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.270000 0.000000 513.410000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.770000 0.000000 508.910000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.265000 0.000000 504.405000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.765000 0.000000 499.905000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.260000 0.000000 495.400000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.755000 0.000000 490.895000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.255000 0.000000 486.395000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.750000 0.000000 481.890000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.250000 0.000000 477.390000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.515000 0.000000 1625.655000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.010000 0.000000 1621.150000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.505000 0.000000 1616.645000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.005000 0.000000 1612.145000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.500000 0.000000 1607.640000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.000000 0.000000 1603.140000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.495000 0.000000 1598.635000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.990000 0.000000 1594.130000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.490000 0.000000 1589.630000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.985000 0.000000 1585.125000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.485000 0.000000 1580.625000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.980000 0.000000 1576.120000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.475000 0.000000 1571.615000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.975000 0.000000 1567.115000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.470000 0.000000 1562.610000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.970000 0.000000 1558.110000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.465000 0.000000 1553.605000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.960000 0.000000 1549.100000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.460000 0.000000 1544.600000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.955000 0.000000 1540.095000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.455000 0.000000 1535.595000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.950000 0.000000 1531.090000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.445000 0.000000 1526.585000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.945000 0.000000 1522.085000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.440000 0.000000 1517.580000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.940000 0.000000 1513.080000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.435000 0.000000 1508.575000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.930000 0.000000 1504.070000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.430000 0.000000 1499.570000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.925000 0.000000 1495.065000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.425000 0.000000 1490.565000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.920000 0.000000 1486.060000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.415000 0.000000 1481.555000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.915000 0.000000 1477.055000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.410000 0.000000 1472.550000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.910000 0.000000 1468.050000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.405000 0.000000 1463.545000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.900000 0.000000 1459.040000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.400000 0.000000 1454.540000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.895000 0.000000 1450.035000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.395000 0.000000 1445.535000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.890000 0.000000 1441.030000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.385000 0.000000 1436.525000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.885000 0.000000 1432.025000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.380000 0.000000 1427.520000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.880000 0.000000 1423.020000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.375000 0.000000 1418.515000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.870000 0.000000 1414.010000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.370000 0.000000 1409.510000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.865000 0.000000 1405.005000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.365000 0.000000 1400.505000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.860000 0.000000 1396.000000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.355000 0.000000 1391.495000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.855000 0.000000 1386.995000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.350000 0.000000 1382.490000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.850000 0.000000 1377.990000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.345000 0.000000 1373.485000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.840000 0.000000 1368.980000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.340000 0.000000 1364.480000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.835000 0.000000 1359.975000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.335000 0.000000 1355.475000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.830000 0.000000 1350.970000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.325000 0.000000 1346.465000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.825000 0.000000 1341.965000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.320000 0.000000 1337.460000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.820000 0.000000 1332.960000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.315000 0.000000 1328.455000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.810000 0.000000 1323.950000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.310000 0.000000 1319.450000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.805000 0.000000 1314.945000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.305000 0.000000 1310.445000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.800000 0.000000 1305.940000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.295000 0.000000 1301.435000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.795000 0.000000 1296.935000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1292.290000 0.000000 1292.430000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.790000 0.000000 1287.930000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.285000 0.000000 1283.425000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.780000 0.000000 1278.920000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.280000 0.000000 1274.420000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.775000 0.000000 1269.915000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.275000 0.000000 1265.415000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.770000 0.000000 1260.910000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.265000 0.000000 1256.405000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.765000 0.000000 1251.905000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.260000 0.000000 1247.400000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.760000 0.000000 1242.900000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.255000 0.000000 1238.395000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.750000 0.000000 1233.890000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.250000 0.000000 1229.390000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.745000 0.000000 1224.885000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.245000 0.000000 1220.385000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.740000 0.000000 1215.880000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.235000 0.000000 1211.375000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.735000 0.000000 1206.875000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.230000 0.000000 1202.370000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.730000 0.000000 1197.870000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.225000 0.000000 1193.365000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.720000 0.000000 1188.860000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.220000 0.000000 1184.360000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.715000 0.000000 1179.855000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.215000 0.000000 1175.355000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.710000 0.000000 1170.850000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.205000 0.000000 1166.345000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.705000 0.000000 1161.845000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.200000 0.000000 1157.340000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.700000 0.000000 1152.840000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.195000 0.000000 1148.335000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.690000 0.000000 1143.830000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.190000 0.000000 1139.330000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.685000 0.000000 1134.825000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.185000 0.000000 1130.325000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.680000 0.000000 1125.820000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.175000 0.000000 1121.315000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.675000 0.000000 1116.815000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.170000 0.000000 1112.310000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.670000 0.000000 1107.810000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.165000 0.000000 1103.305000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.660000 0.000000 1098.800000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.160000 0.000000 1094.300000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.655000 0.000000 1089.795000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.155000 0.000000 1085.295000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.650000 0.000000 1080.790000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.145000 0.000000 1076.285000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.645000 0.000000 1071.785000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.140000 0.000000 1067.280000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.640000 0.000000 1062.780000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.135000 0.000000 1058.275000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.630000 0.000000 1053.770000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.895000 0.000000 2202.035000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2197.395000 0.000000 2197.535000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2192.890000 0.000000 2193.030000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.390000 0.000000 2188.530000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.885000 0.000000 2184.025000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.380000 0.000000 2179.520000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2174.880000 0.000000 2175.020000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.375000 0.000000 2170.515000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.875000 0.000000 2166.015000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.370000 0.000000 2161.510000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.865000 0.000000 2157.005000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.365000 0.000000 2152.505000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.860000 0.000000 2148.000000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.360000 0.000000 2143.500000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.855000 0.000000 2138.995000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.350000 0.000000 2134.490000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.850000 0.000000 2129.990000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.345000 0.000000 2125.485000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2120.845000 0.000000 2120.985000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2116.340000 0.000000 2116.480000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2111.835000 0.000000 2111.975000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.335000 0.000000 2107.475000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.830000 0.000000 2102.970000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2098.330000 0.000000 2098.470000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.825000 0.000000 2093.965000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.320000 0.000000 2089.460000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.820000 0.000000 2084.960000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.315000 0.000000 2080.455000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.815000 0.000000 2075.955000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.310000 0.000000 2071.450000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.805000 0.000000 2066.945000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2062.305000 0.000000 2062.445000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.800000 0.000000 2057.940000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.300000 0.000000 2053.440000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.795000 0.000000 2048.935000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.290000 0.000000 2044.430000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.790000 0.000000 2039.930000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.285000 0.000000 2035.425000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.785000 0.000000 2030.925000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.280000 0.000000 2026.420000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.775000 0.000000 2021.915000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.275000 0.000000 2017.415000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.770000 0.000000 2012.910000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.270000 0.000000 2008.410000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.765000 0.000000 2003.905000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.260000 0.000000 1999.400000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.760000 0.000000 1994.900000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.255000 0.000000 1990.395000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.755000 0.000000 1985.895000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.250000 0.000000 1981.390000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.745000 0.000000 1976.885000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.245000 0.000000 1972.385000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.740000 0.000000 1967.880000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.240000 0.000000 1963.380000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.735000 0.000000 1958.875000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.230000 0.000000 1954.370000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.730000 0.000000 1949.870000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.225000 0.000000 1945.365000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.725000 0.000000 1940.865000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.220000 0.000000 1936.360000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.715000 0.000000 1931.855000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.215000 0.000000 1927.355000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.710000 0.000000 1922.850000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1918.210000 0.000000 1918.350000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.705000 0.000000 1913.845000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.200000 0.000000 1909.340000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.700000 0.000000 1904.840000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.195000 0.000000 1900.335000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1895.695000 0.000000 1895.835000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.190000 0.000000 1891.330000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.685000 0.000000 1886.825000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.185000 0.000000 1882.325000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.680000 0.000000 1877.820000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.180000 0.000000 1873.320000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.675000 0.000000 1868.815000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.170000 0.000000 1864.310000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.670000 0.000000 1859.810000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.165000 0.000000 1855.305000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.665000 0.000000 1850.805000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.160000 0.000000 1846.300000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.655000 0.000000 1841.795000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.155000 0.000000 1837.295000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.650000 0.000000 1832.790000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.150000 0.000000 1828.290000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.645000 0.000000 1823.785000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.140000 0.000000 1819.280000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1814.640000 0.000000 1814.780000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.135000 0.000000 1810.275000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.635000 0.000000 1805.775000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.130000 0.000000 1801.270000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.625000 0.000000 1796.765000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.125000 0.000000 1792.265000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.620000 0.000000 1787.760000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.120000 0.000000 1783.260000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1778.615000 0.000000 1778.755000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.110000 0.000000 1774.250000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.610000 0.000000 1769.750000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.105000 0.000000 1765.245000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.605000 0.000000 1760.745000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.100000 0.000000 1756.240000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.595000 0.000000 1751.735000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.095000 0.000000 1747.235000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.590000 0.000000 1742.730000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.090000 0.000000 1738.230000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.585000 0.000000 1733.725000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.080000 0.000000 1729.220000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.580000 0.000000 1724.720000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.075000 0.000000 1720.215000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.575000 0.000000 1715.715000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.070000 0.000000 1711.210000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.565000 0.000000 1706.705000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.065000 0.000000 1702.205000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.560000 0.000000 1697.700000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.060000 0.000000 1693.200000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.555000 0.000000 1688.695000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.050000 0.000000 1684.190000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.550000 0.000000 1679.690000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.045000 0.000000 1675.185000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.545000 0.000000 1670.685000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.040000 0.000000 1666.180000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.535000 0.000000 1661.675000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.035000 0.000000 1657.175000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.530000 0.000000 1652.670000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.030000 0.000000 1648.170000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.525000 0.000000 1643.665000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.020000 0.000000 1639.160000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.520000 0.000000 1634.660000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.015000 0.000000 1630.155000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 110.780000 0.800000 111.080000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 277.170000 0.800000 277.470000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 443.560000 0.800000 443.860000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 665.420000 0.800000 665.720000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 887.275000 0.800000 887.575000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1109.130000 0.800000 1109.430000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1330.985000 0.800000 1331.285000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1552.840000 0.800000 1553.140000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1774.700000 0.800000 1775.000000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1996.555000 0.800000 1996.855000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2218.410000 0.800000 2218.710000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2440.265000 0.800000 2440.565000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2662.120000 0.800000 2662.420000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2883.980000 0.800000 2884.280000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.810000 2939.150000 126.950000 2939.640000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.570000 2939.150000 380.710000 2939.640000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.330000 2939.150000 634.470000 2939.640000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.090000 2939.150000 888.230000 2939.640000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.850000 2939.150000 1141.990000 2939.640000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.610000 2939.150000 1395.750000 2939.640000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.370000 2939.150000 1649.510000 2939.640000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.130000 2939.150000 1903.270000 2939.640000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.890000 2939.150000 2157.030000 2939.640000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2826.400000 2220.420000 2826.700000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2600.275000 2220.420000 2600.575000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2374.150000 2220.420000 2374.450000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2148.030000 2220.420000 2148.330000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1921.905000 2220.420000 1922.205000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1695.780000 2220.420000 1696.080000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1469.655000 2220.420000 1469.955000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1243.530000 2220.420000 1243.830000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1017.410000 2220.420000 1017.710000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 847.815000 2220.420000 848.115000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 678.220000 2220.420000 678.520000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 508.630000 2220.420000 508.930000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 339.035000 2220.420000 339.335000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 169.445000 2220.420000 169.745000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2.560000 2220.420000 2.860000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 55.315000 0.800000 55.615000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 221.705000 0.800000 222.005000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 388.100000 0.800000 388.400000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 609.955000 0.800000 610.255000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 831.810000 0.800000 832.110000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1053.665000 0.800000 1053.965000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1275.520000 0.800000 1275.820000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1497.380000 0.800000 1497.680000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1719.235000 0.800000 1719.535000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1941.090000 0.800000 1941.390000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2162.945000 0.800000 2163.245000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2384.800000 0.800000 2385.100000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2606.660000 0.800000 2606.960000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2828.515000 0.800000 2828.815000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.370000 2939.150000 63.510000 2939.640000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.130000 2939.150000 317.270000 2939.640000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.890000 2939.150000 571.030000 2939.640000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.650000 2939.150000 824.790000 2939.640000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.410000 2939.150000 1078.550000 2939.640000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.170000 2939.150000 1332.310000 2939.640000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.930000 2939.150000 1586.070000 2939.640000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.690000 2939.150000 1839.830000 2939.640000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.450000 2939.150000 2093.590000 2939.640000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2882.930000 2220.420000 2883.230000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2656.805000 2220.420000 2657.105000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2430.685000 2220.420000 2430.985000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2204.560000 2220.420000 2204.860000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1978.435000 2220.420000 1978.735000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1752.310000 2220.420000 1752.610000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1526.185000 2220.420000 1526.485000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1300.065000 2220.420000 1300.365000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1073.940000 2220.420000 1074.240000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 904.345000 2220.420000 904.645000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 734.755000 2220.420000 735.055000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 565.160000 2220.420000 565.460000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 395.565000 2220.420000 395.865000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 225.975000 2220.420000 226.275000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 56.380000 2220.420000 56.680000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 3.170000 0.800000 3.470000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 166.240000 0.800000 166.540000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 332.635000 0.800000 332.935000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 554.490000 0.800000 554.790000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 776.345000 0.800000 776.645000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 998.200000 0.800000 998.500000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1220.060000 0.800000 1220.360000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1441.915000 0.800000 1442.215000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1663.770000 0.800000 1664.070000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1885.625000 0.800000 1885.925000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2107.480000 0.800000 2107.780000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2329.340000 0.800000 2329.640000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2551.195000 0.800000 2551.495000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2773.050000 0.800000 2773.350000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.380000 2939.150000 3.520000 2939.640000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.690000 2939.150000 253.830000 2939.640000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.450000 2939.150000 507.590000 2939.640000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.210000 2939.150000 761.350000 2939.640000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.970000 2939.150000 1015.110000 2939.640000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.730000 2939.150000 1268.870000 2939.640000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.490000 2939.150000 1522.630000 2939.640000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.250000 2939.150000 1776.390000 2939.640000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.010000 2939.150000 2030.150000 2939.640000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2934.830000 2220.420000 2935.130000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2713.340000 2220.420000 2713.640000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2487.215000 2220.420000 2487.515000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2261.090000 2220.420000 2261.390000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2034.965000 2220.420000 2035.265000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1808.840000 2220.420000 1809.140000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1582.720000 2220.420000 1583.020000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1356.595000 2220.420000 1356.895000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1130.470000 2220.420000 1130.770000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 960.875000 2220.420000 961.175000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 791.285000 2220.420000 791.585000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 621.690000 2220.420000 621.990000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 452.100000 2220.420000 452.400000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 282.505000 2220.420000 282.805000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 112.910000 2220.420000 113.210000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 499.025000 0.800000 499.325000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 720.880000 0.800000 721.180000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 942.740000 0.800000 943.040000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1164.595000 0.800000 1164.895000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1386.450000 0.800000 1386.750000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1608.305000 0.800000 1608.605000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1830.160000 0.800000 1830.460000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2052.020000 0.800000 2052.320000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2273.875000 0.800000 2274.175000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2495.730000 0.800000 2496.030000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2717.585000 0.800000 2717.885000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2935.440000 0.800000 2935.740000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.250000 2939.150000 190.390000 2939.640000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.010000 2939.150000 444.150000 2939.640000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.770000 2939.150000 697.910000 2939.640000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.530000 2939.150000 951.670000 2939.640000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.290000 2939.150000 1205.430000 2939.640000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.050000 2939.150000 1459.190000 2939.640000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.810000 2939.150000 1712.950000 2939.640000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.570000 2939.150000 1966.710000 2939.640000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.980000 2939.150000 2216.120000 2939.640000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2769.870000 2220.420000 2770.170000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2543.745000 2220.420000 2544.045000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2317.620000 2220.420000 2317.920000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 2091.495000 2220.420000 2091.795000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1865.375000 2220.420000 1865.675000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1639.250000 2220.420000 1639.550000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1413.125000 2220.420000 1413.425000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2219.620000 1187.000000 2220.420000 1187.300000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.400000 0.000000 2206.540000 0.490000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.060000 0.000000 2215.200000 0.490000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.405000 0.000000 2215.545000 0.490000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2210.905000 0.000000 2211.045000 0.490000 ;
    END
  END user_irq[0]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2212.360000 5.930000 2214.360000 2933.030000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.060000 5.930000 8.060000 2933.030000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1675.210000 1021.045000 1676.950000 1409.025000 ;
      LAYER met4 ;
        RECT 2143.730000 1021.045000 2145.470000 1409.025000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 535.980000 2470.465000 537.720000 2858.445000 ;
      LAYER met4 ;
        RECT 67.460000 2470.465000 69.200000 2858.445000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2146.210000 534.690000 2147.950000 922.670000 ;
      LAYER met4 ;
        RECT 1677.690000 534.690000 1679.430000 922.670000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2141.480000 1507.405000 2143.220000 1895.385000 ;
      LAYER met4 ;
        RECT 1672.960000 1507.405000 1674.700000 1895.385000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2152.840000 2469.100000 2154.580000 2857.080000 ;
      LAYER met4 ;
        RECT 1684.320000 2469.100000 1686.060000 2857.080000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1662.065000 1970.370000 1663.805000 2358.350000 ;
      LAYER met4 ;
        RECT 2130.585000 1970.370000 2132.325000 2358.350000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1083.330000 2463.890000 1085.070000 2851.870000 ;
      LAYER met4 ;
        RECT 614.810000 2463.890000 616.550000 2851.870000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1149.420000 2464.745000 1151.160000 2852.725000 ;
      LAYER met4 ;
        RECT 1617.940000 2464.745000 1619.680000 2852.725000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2.060000 1.930000 4.060000 2937.030000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.360000 1.930000 2218.360000 2937.030000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2147.130000 1017.645000 2148.870000 1412.425000 ;
      LAYER met4 ;
        RECT 1671.810000 1017.645000 1673.550000 1412.425000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 64.060000 2467.065000 65.800000 2861.845000 ;
      LAYER met4 ;
        RECT 539.380000 2467.065000 541.120000 2861.845000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1674.290000 531.290000 1676.030000 926.070000 ;
      LAYER met4 ;
        RECT 2149.610000 531.290000 2151.350000 926.070000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1669.560000 1504.005000 1671.300000 1898.785000 ;
      LAYER met4 ;
        RECT 2144.880000 1504.005000 2146.620000 1898.785000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1680.920000 2465.700000 1682.660000 2860.480000 ;
      LAYER met4 ;
        RECT 2156.240000 2465.700000 2157.980000 2860.480000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2133.985000 1966.970000 2135.725000 2361.750000 ;
      LAYER met4 ;
        RECT 1658.665000 1966.970000 1660.405000 2361.750000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 611.410000 2460.490000 613.150000 2855.270000 ;
      LAYER met4 ;
        RECT 1086.730000 2460.490000 1088.470000 2855.270000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1621.340000 2461.345000 1623.080000 2856.125000 ;
      LAYER met4 ;
        RECT 1146.020000 2461.345000 1147.760000 2856.125000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END VGND
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2220.420000 2939.640000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2220.420000 2939.640000 ;
    LAYER met2 ;
      RECT 2216.260000 2939.010000 2220.420000 2939.640000 ;
      RECT 2157.170000 2939.010000 2215.840000 2939.640000 ;
      RECT 2093.730000 2939.010000 2156.750000 2939.640000 ;
      RECT 2030.290000 2939.010000 2093.310000 2939.640000 ;
      RECT 1966.850000 2939.010000 2029.870000 2939.640000 ;
      RECT 1903.410000 2939.010000 1966.430000 2939.640000 ;
      RECT 1839.970000 2939.010000 1902.990000 2939.640000 ;
      RECT 1776.530000 2939.010000 1839.550000 2939.640000 ;
      RECT 1713.090000 2939.010000 1776.110000 2939.640000 ;
      RECT 1649.650000 2939.010000 1712.670000 2939.640000 ;
      RECT 1586.210000 2939.010000 1649.230000 2939.640000 ;
      RECT 1522.770000 2939.010000 1585.790000 2939.640000 ;
      RECT 1459.330000 2939.010000 1522.350000 2939.640000 ;
      RECT 1395.890000 2939.010000 1458.910000 2939.640000 ;
      RECT 1332.450000 2939.010000 1395.470000 2939.640000 ;
      RECT 1269.010000 2939.010000 1332.030000 2939.640000 ;
      RECT 1205.570000 2939.010000 1268.590000 2939.640000 ;
      RECT 1142.130000 2939.010000 1205.150000 2939.640000 ;
      RECT 1078.690000 2939.010000 1141.710000 2939.640000 ;
      RECT 1015.250000 2939.010000 1078.270000 2939.640000 ;
      RECT 951.810000 2939.010000 1014.830000 2939.640000 ;
      RECT 888.370000 2939.010000 951.390000 2939.640000 ;
      RECT 824.930000 2939.010000 887.950000 2939.640000 ;
      RECT 761.490000 2939.010000 824.510000 2939.640000 ;
      RECT 698.050000 2939.010000 761.070000 2939.640000 ;
      RECT 634.610000 2939.010000 697.630000 2939.640000 ;
      RECT 571.170000 2939.010000 634.190000 2939.640000 ;
      RECT 507.730000 2939.010000 570.750000 2939.640000 ;
      RECT 444.290000 2939.010000 507.310000 2939.640000 ;
      RECT 380.850000 2939.010000 443.870000 2939.640000 ;
      RECT 317.410000 2939.010000 380.430000 2939.640000 ;
      RECT 253.970000 2939.010000 316.990000 2939.640000 ;
      RECT 190.530000 2939.010000 253.550000 2939.640000 ;
      RECT 127.090000 2939.010000 190.110000 2939.640000 ;
      RECT 63.650000 2939.010000 126.670000 2939.640000 ;
      RECT 3.660000 2939.010000 63.230000 2939.640000 ;
      RECT 0.000000 2939.010000 3.240000 2939.640000 ;
      RECT 0.000000 0.630000 2220.420000 2939.010000 ;
      RECT 2215.685000 0.000000 2220.420000 0.630000 ;
      RECT 2211.185000 0.000000 2214.920000 0.630000 ;
      RECT 2206.680000 0.000000 2210.765000 0.630000 ;
      RECT 2202.175000 0.000000 2206.260000 0.630000 ;
      RECT 2197.675000 0.000000 2201.755000 0.630000 ;
      RECT 2193.170000 0.000000 2197.255000 0.630000 ;
      RECT 2188.670000 0.000000 2192.750000 0.630000 ;
      RECT 2184.165000 0.000000 2188.250000 0.630000 ;
      RECT 2179.660000 0.000000 2183.745000 0.630000 ;
      RECT 2175.160000 0.000000 2179.240000 0.630000 ;
      RECT 2170.655000 0.000000 2174.740000 0.630000 ;
      RECT 2166.155000 0.000000 2170.235000 0.630000 ;
      RECT 2161.650000 0.000000 2165.735000 0.630000 ;
      RECT 2157.145000 0.000000 2161.230000 0.630000 ;
      RECT 2152.645000 0.000000 2156.725000 0.630000 ;
      RECT 2148.140000 0.000000 2152.225000 0.630000 ;
      RECT 2143.640000 0.000000 2147.720000 0.630000 ;
      RECT 2139.135000 0.000000 2143.220000 0.630000 ;
      RECT 2134.630000 0.000000 2138.715000 0.630000 ;
      RECT 2130.130000 0.000000 2134.210000 0.630000 ;
      RECT 2125.625000 0.000000 2129.710000 0.630000 ;
      RECT 2121.125000 0.000000 2125.205000 0.630000 ;
      RECT 2116.620000 0.000000 2120.705000 0.630000 ;
      RECT 2112.115000 0.000000 2116.200000 0.630000 ;
      RECT 2107.615000 0.000000 2111.695000 0.630000 ;
      RECT 2103.110000 0.000000 2107.195000 0.630000 ;
      RECT 2098.610000 0.000000 2102.690000 0.630000 ;
      RECT 2094.105000 0.000000 2098.190000 0.630000 ;
      RECT 2089.600000 0.000000 2093.685000 0.630000 ;
      RECT 2085.100000 0.000000 2089.180000 0.630000 ;
      RECT 2080.595000 0.000000 2084.680000 0.630000 ;
      RECT 2076.095000 0.000000 2080.175000 0.630000 ;
      RECT 2071.590000 0.000000 2075.675000 0.630000 ;
      RECT 2067.085000 0.000000 2071.170000 0.630000 ;
      RECT 2062.585000 0.000000 2066.665000 0.630000 ;
      RECT 2058.080000 0.000000 2062.165000 0.630000 ;
      RECT 2053.580000 0.000000 2057.660000 0.630000 ;
      RECT 2049.075000 0.000000 2053.160000 0.630000 ;
      RECT 2044.570000 0.000000 2048.655000 0.630000 ;
      RECT 2040.070000 0.000000 2044.150000 0.630000 ;
      RECT 2035.565000 0.000000 2039.650000 0.630000 ;
      RECT 2031.065000 0.000000 2035.145000 0.630000 ;
      RECT 2026.560000 0.000000 2030.645000 0.630000 ;
      RECT 2022.055000 0.000000 2026.140000 0.630000 ;
      RECT 2017.555000 0.000000 2021.635000 0.630000 ;
      RECT 2013.050000 0.000000 2017.135000 0.630000 ;
      RECT 2008.550000 0.000000 2012.630000 0.630000 ;
      RECT 2004.045000 0.000000 2008.130000 0.630000 ;
      RECT 1999.540000 0.000000 2003.625000 0.630000 ;
      RECT 1995.040000 0.000000 1999.120000 0.630000 ;
      RECT 1990.535000 0.000000 1994.620000 0.630000 ;
      RECT 1986.035000 0.000000 1990.115000 0.630000 ;
      RECT 1981.530000 0.000000 1985.615000 0.630000 ;
      RECT 1977.025000 0.000000 1981.110000 0.630000 ;
      RECT 1972.525000 0.000000 1976.605000 0.630000 ;
      RECT 1968.020000 0.000000 1972.105000 0.630000 ;
      RECT 1963.520000 0.000000 1967.600000 0.630000 ;
      RECT 1959.015000 0.000000 1963.100000 0.630000 ;
      RECT 1954.510000 0.000000 1958.595000 0.630000 ;
      RECT 1950.010000 0.000000 1954.090000 0.630000 ;
      RECT 1945.505000 0.000000 1949.590000 0.630000 ;
      RECT 1941.005000 0.000000 1945.085000 0.630000 ;
      RECT 1936.500000 0.000000 1940.585000 0.630000 ;
      RECT 1931.995000 0.000000 1936.080000 0.630000 ;
      RECT 1927.495000 0.000000 1931.575000 0.630000 ;
      RECT 1922.990000 0.000000 1927.075000 0.630000 ;
      RECT 1918.490000 0.000000 1922.570000 0.630000 ;
      RECT 1913.985000 0.000000 1918.070000 0.630000 ;
      RECT 1909.480000 0.000000 1913.565000 0.630000 ;
      RECT 1904.980000 0.000000 1909.060000 0.630000 ;
      RECT 1900.475000 0.000000 1904.560000 0.630000 ;
      RECT 1895.975000 0.000000 1900.055000 0.630000 ;
      RECT 1891.470000 0.000000 1895.555000 0.630000 ;
      RECT 1886.965000 0.000000 1891.050000 0.630000 ;
      RECT 1882.465000 0.000000 1886.545000 0.630000 ;
      RECT 1877.960000 0.000000 1882.045000 0.630000 ;
      RECT 1873.460000 0.000000 1877.540000 0.630000 ;
      RECT 1868.955000 0.000000 1873.040000 0.630000 ;
      RECT 1864.450000 0.000000 1868.535000 0.630000 ;
      RECT 1859.950000 0.000000 1864.030000 0.630000 ;
      RECT 1855.445000 0.000000 1859.530000 0.630000 ;
      RECT 1850.945000 0.000000 1855.025000 0.630000 ;
      RECT 1846.440000 0.000000 1850.525000 0.630000 ;
      RECT 1841.935000 0.000000 1846.020000 0.630000 ;
      RECT 1837.435000 0.000000 1841.515000 0.630000 ;
      RECT 1832.930000 0.000000 1837.015000 0.630000 ;
      RECT 1828.430000 0.000000 1832.510000 0.630000 ;
      RECT 1823.925000 0.000000 1828.010000 0.630000 ;
      RECT 1819.420000 0.000000 1823.505000 0.630000 ;
      RECT 1814.920000 0.000000 1819.000000 0.630000 ;
      RECT 1810.415000 0.000000 1814.500000 0.630000 ;
      RECT 1805.915000 0.000000 1809.995000 0.630000 ;
      RECT 1801.410000 0.000000 1805.495000 0.630000 ;
      RECT 1796.905000 0.000000 1800.990000 0.630000 ;
      RECT 1792.405000 0.000000 1796.485000 0.630000 ;
      RECT 1787.900000 0.000000 1791.985000 0.630000 ;
      RECT 1783.400000 0.000000 1787.480000 0.630000 ;
      RECT 1778.895000 0.000000 1782.980000 0.630000 ;
      RECT 1774.390000 0.000000 1778.475000 0.630000 ;
      RECT 1769.890000 0.000000 1773.970000 0.630000 ;
      RECT 1765.385000 0.000000 1769.470000 0.630000 ;
      RECT 1760.885000 0.000000 1764.965000 0.630000 ;
      RECT 1756.380000 0.000000 1760.465000 0.630000 ;
      RECT 1751.875000 0.000000 1755.960000 0.630000 ;
      RECT 1747.375000 0.000000 1751.455000 0.630000 ;
      RECT 1742.870000 0.000000 1746.955000 0.630000 ;
      RECT 1738.370000 0.000000 1742.450000 0.630000 ;
      RECT 1733.865000 0.000000 1737.950000 0.630000 ;
      RECT 1729.360000 0.000000 1733.445000 0.630000 ;
      RECT 1724.860000 0.000000 1728.940000 0.630000 ;
      RECT 1720.355000 0.000000 1724.440000 0.630000 ;
      RECT 1715.855000 0.000000 1719.935000 0.630000 ;
      RECT 1711.350000 0.000000 1715.435000 0.630000 ;
      RECT 1706.845000 0.000000 1710.930000 0.630000 ;
      RECT 1702.345000 0.000000 1706.425000 0.630000 ;
      RECT 1697.840000 0.000000 1701.925000 0.630000 ;
      RECT 1693.340000 0.000000 1697.420000 0.630000 ;
      RECT 1688.835000 0.000000 1692.920000 0.630000 ;
      RECT 1684.330000 0.000000 1688.415000 0.630000 ;
      RECT 1679.830000 0.000000 1683.910000 0.630000 ;
      RECT 1675.325000 0.000000 1679.410000 0.630000 ;
      RECT 1670.825000 0.000000 1674.905000 0.630000 ;
      RECT 1666.320000 0.000000 1670.405000 0.630000 ;
      RECT 1661.815000 0.000000 1665.900000 0.630000 ;
      RECT 1657.315000 0.000000 1661.395000 0.630000 ;
      RECT 1652.810000 0.000000 1656.895000 0.630000 ;
      RECT 1648.310000 0.000000 1652.390000 0.630000 ;
      RECT 1643.805000 0.000000 1647.890000 0.630000 ;
      RECT 1639.300000 0.000000 1643.385000 0.630000 ;
      RECT 1634.800000 0.000000 1638.880000 0.630000 ;
      RECT 1630.295000 0.000000 1634.380000 0.630000 ;
      RECT 1625.795000 0.000000 1629.875000 0.630000 ;
      RECT 1621.290000 0.000000 1625.375000 0.630000 ;
      RECT 1616.785000 0.000000 1620.870000 0.630000 ;
      RECT 1612.285000 0.000000 1616.365000 0.630000 ;
      RECT 1607.780000 0.000000 1611.865000 0.630000 ;
      RECT 1603.280000 0.000000 1607.360000 0.630000 ;
      RECT 1598.775000 0.000000 1602.860000 0.630000 ;
      RECT 1594.270000 0.000000 1598.355000 0.630000 ;
      RECT 1589.770000 0.000000 1593.850000 0.630000 ;
      RECT 1585.265000 0.000000 1589.350000 0.630000 ;
      RECT 1580.765000 0.000000 1584.845000 0.630000 ;
      RECT 1576.260000 0.000000 1580.345000 0.630000 ;
      RECT 1571.755000 0.000000 1575.840000 0.630000 ;
      RECT 1567.255000 0.000000 1571.335000 0.630000 ;
      RECT 1562.750000 0.000000 1566.835000 0.630000 ;
      RECT 1558.250000 0.000000 1562.330000 0.630000 ;
      RECT 1553.745000 0.000000 1557.830000 0.630000 ;
      RECT 1549.240000 0.000000 1553.325000 0.630000 ;
      RECT 1544.740000 0.000000 1548.820000 0.630000 ;
      RECT 1540.235000 0.000000 1544.320000 0.630000 ;
      RECT 1535.735000 0.000000 1539.815000 0.630000 ;
      RECT 1531.230000 0.000000 1535.315000 0.630000 ;
      RECT 1526.725000 0.000000 1530.810000 0.630000 ;
      RECT 1522.225000 0.000000 1526.305000 0.630000 ;
      RECT 1517.720000 0.000000 1521.805000 0.630000 ;
      RECT 1513.220000 0.000000 1517.300000 0.630000 ;
      RECT 1508.715000 0.000000 1512.800000 0.630000 ;
      RECT 1504.210000 0.000000 1508.295000 0.630000 ;
      RECT 1499.710000 0.000000 1503.790000 0.630000 ;
      RECT 1495.205000 0.000000 1499.290000 0.630000 ;
      RECT 1490.705000 0.000000 1494.785000 0.630000 ;
      RECT 1486.200000 0.000000 1490.285000 0.630000 ;
      RECT 1481.695000 0.000000 1485.780000 0.630000 ;
      RECT 1477.195000 0.000000 1481.275000 0.630000 ;
      RECT 1472.690000 0.000000 1476.775000 0.630000 ;
      RECT 1468.190000 0.000000 1472.270000 0.630000 ;
      RECT 1463.685000 0.000000 1467.770000 0.630000 ;
      RECT 1459.180000 0.000000 1463.265000 0.630000 ;
      RECT 1454.680000 0.000000 1458.760000 0.630000 ;
      RECT 1450.175000 0.000000 1454.260000 0.630000 ;
      RECT 1445.675000 0.000000 1449.755000 0.630000 ;
      RECT 1441.170000 0.000000 1445.255000 0.630000 ;
      RECT 1436.665000 0.000000 1440.750000 0.630000 ;
      RECT 1432.165000 0.000000 1436.245000 0.630000 ;
      RECT 1427.660000 0.000000 1431.745000 0.630000 ;
      RECT 1423.160000 0.000000 1427.240000 0.630000 ;
      RECT 1418.655000 0.000000 1422.740000 0.630000 ;
      RECT 1414.150000 0.000000 1418.235000 0.630000 ;
      RECT 1409.650000 0.000000 1413.730000 0.630000 ;
      RECT 1405.145000 0.000000 1409.230000 0.630000 ;
      RECT 1400.645000 0.000000 1404.725000 0.630000 ;
      RECT 1396.140000 0.000000 1400.225000 0.630000 ;
      RECT 1391.635000 0.000000 1395.720000 0.630000 ;
      RECT 1387.135000 0.000000 1391.215000 0.630000 ;
      RECT 1382.630000 0.000000 1386.715000 0.630000 ;
      RECT 1378.130000 0.000000 1382.210000 0.630000 ;
      RECT 1373.625000 0.000000 1377.710000 0.630000 ;
      RECT 1369.120000 0.000000 1373.205000 0.630000 ;
      RECT 1364.620000 0.000000 1368.700000 0.630000 ;
      RECT 1360.115000 0.000000 1364.200000 0.630000 ;
      RECT 1355.615000 0.000000 1359.695000 0.630000 ;
      RECT 1351.110000 0.000000 1355.195000 0.630000 ;
      RECT 1346.605000 0.000000 1350.690000 0.630000 ;
      RECT 1342.105000 0.000000 1346.185000 0.630000 ;
      RECT 1337.600000 0.000000 1341.685000 0.630000 ;
      RECT 1333.100000 0.000000 1337.180000 0.630000 ;
      RECT 1328.595000 0.000000 1332.680000 0.630000 ;
      RECT 1324.090000 0.000000 1328.175000 0.630000 ;
      RECT 1319.590000 0.000000 1323.670000 0.630000 ;
      RECT 1315.085000 0.000000 1319.170000 0.630000 ;
      RECT 1310.585000 0.000000 1314.665000 0.630000 ;
      RECT 1306.080000 0.000000 1310.165000 0.630000 ;
      RECT 1301.575000 0.000000 1305.660000 0.630000 ;
      RECT 1297.075000 0.000000 1301.155000 0.630000 ;
      RECT 1292.570000 0.000000 1296.655000 0.630000 ;
      RECT 1288.070000 0.000000 1292.150000 0.630000 ;
      RECT 1283.565000 0.000000 1287.650000 0.630000 ;
      RECT 1279.060000 0.000000 1283.145000 0.630000 ;
      RECT 1274.560000 0.000000 1278.640000 0.630000 ;
      RECT 1270.055000 0.000000 1274.140000 0.630000 ;
      RECT 1265.555000 0.000000 1269.635000 0.630000 ;
      RECT 1261.050000 0.000000 1265.135000 0.630000 ;
      RECT 1256.545000 0.000000 1260.630000 0.630000 ;
      RECT 1252.045000 0.000000 1256.125000 0.630000 ;
      RECT 1247.540000 0.000000 1251.625000 0.630000 ;
      RECT 1243.040000 0.000000 1247.120000 0.630000 ;
      RECT 1238.535000 0.000000 1242.620000 0.630000 ;
      RECT 1234.030000 0.000000 1238.115000 0.630000 ;
      RECT 1229.530000 0.000000 1233.610000 0.630000 ;
      RECT 1225.025000 0.000000 1229.110000 0.630000 ;
      RECT 1220.525000 0.000000 1224.605000 0.630000 ;
      RECT 1216.020000 0.000000 1220.105000 0.630000 ;
      RECT 1211.515000 0.000000 1215.600000 0.630000 ;
      RECT 1207.015000 0.000000 1211.095000 0.630000 ;
      RECT 1202.510000 0.000000 1206.595000 0.630000 ;
      RECT 1198.010000 0.000000 1202.090000 0.630000 ;
      RECT 1193.505000 0.000000 1197.590000 0.630000 ;
      RECT 1189.000000 0.000000 1193.085000 0.630000 ;
      RECT 1184.500000 0.000000 1188.580000 0.630000 ;
      RECT 1179.995000 0.000000 1184.080000 0.630000 ;
      RECT 1175.495000 0.000000 1179.575000 0.630000 ;
      RECT 1170.990000 0.000000 1175.075000 0.630000 ;
      RECT 1166.485000 0.000000 1170.570000 0.630000 ;
      RECT 1161.985000 0.000000 1166.065000 0.630000 ;
      RECT 1157.480000 0.000000 1161.565000 0.630000 ;
      RECT 1152.980000 0.000000 1157.060000 0.630000 ;
      RECT 1148.475000 0.000000 1152.560000 0.630000 ;
      RECT 1143.970000 0.000000 1148.055000 0.630000 ;
      RECT 1139.470000 0.000000 1143.550000 0.630000 ;
      RECT 1134.965000 0.000000 1139.050000 0.630000 ;
      RECT 1130.465000 0.000000 1134.545000 0.630000 ;
      RECT 1125.960000 0.000000 1130.045000 0.630000 ;
      RECT 1121.455000 0.000000 1125.540000 0.630000 ;
      RECT 1116.955000 0.000000 1121.035000 0.630000 ;
      RECT 1112.450000 0.000000 1116.535000 0.630000 ;
      RECT 1107.950000 0.000000 1112.030000 0.630000 ;
      RECT 1103.445000 0.000000 1107.530000 0.630000 ;
      RECT 1098.940000 0.000000 1103.025000 0.630000 ;
      RECT 1094.440000 0.000000 1098.520000 0.630000 ;
      RECT 1089.935000 0.000000 1094.020000 0.630000 ;
      RECT 1085.435000 0.000000 1089.515000 0.630000 ;
      RECT 1080.930000 0.000000 1085.015000 0.630000 ;
      RECT 1076.425000 0.000000 1080.510000 0.630000 ;
      RECT 1071.925000 0.000000 1076.005000 0.630000 ;
      RECT 1067.420000 0.000000 1071.505000 0.630000 ;
      RECT 1062.920000 0.000000 1067.000000 0.630000 ;
      RECT 1058.415000 0.000000 1062.500000 0.630000 ;
      RECT 1053.910000 0.000000 1057.995000 0.630000 ;
      RECT 1049.410000 0.000000 1053.490000 0.630000 ;
      RECT 1044.905000 0.000000 1048.990000 0.630000 ;
      RECT 1040.405000 0.000000 1044.485000 0.630000 ;
      RECT 1035.900000 0.000000 1039.985000 0.630000 ;
      RECT 1031.395000 0.000000 1035.480000 0.630000 ;
      RECT 1026.895000 0.000000 1030.975000 0.630000 ;
      RECT 1022.390000 0.000000 1026.475000 0.630000 ;
      RECT 1017.890000 0.000000 1021.970000 0.630000 ;
      RECT 1013.385000 0.000000 1017.470000 0.630000 ;
      RECT 1008.880000 0.000000 1012.965000 0.630000 ;
      RECT 1004.380000 0.000000 1008.460000 0.630000 ;
      RECT 999.875000 0.000000 1003.960000 0.630000 ;
      RECT 995.375000 0.000000 999.455000 0.630000 ;
      RECT 990.870000 0.000000 994.955000 0.630000 ;
      RECT 986.365000 0.000000 990.450000 0.630000 ;
      RECT 981.865000 0.000000 985.945000 0.630000 ;
      RECT 977.360000 0.000000 981.445000 0.630000 ;
      RECT 972.860000 0.000000 976.940000 0.630000 ;
      RECT 968.355000 0.000000 972.440000 0.630000 ;
      RECT 963.850000 0.000000 967.935000 0.630000 ;
      RECT 959.350000 0.000000 963.430000 0.630000 ;
      RECT 954.845000 0.000000 958.930000 0.630000 ;
      RECT 950.345000 0.000000 954.425000 0.630000 ;
      RECT 945.840000 0.000000 949.925000 0.630000 ;
      RECT 941.335000 0.000000 945.420000 0.630000 ;
      RECT 936.835000 0.000000 940.915000 0.630000 ;
      RECT 932.330000 0.000000 936.415000 0.630000 ;
      RECT 927.830000 0.000000 931.910000 0.630000 ;
      RECT 923.325000 0.000000 927.410000 0.630000 ;
      RECT 918.820000 0.000000 922.905000 0.630000 ;
      RECT 914.320000 0.000000 918.400000 0.630000 ;
      RECT 909.815000 0.000000 913.900000 0.630000 ;
      RECT 905.315000 0.000000 909.395000 0.630000 ;
      RECT 900.810000 0.000000 904.895000 0.630000 ;
      RECT 896.305000 0.000000 900.390000 0.630000 ;
      RECT 891.805000 0.000000 895.885000 0.630000 ;
      RECT 887.300000 0.000000 891.385000 0.630000 ;
      RECT 882.800000 0.000000 886.880000 0.630000 ;
      RECT 878.295000 0.000000 882.380000 0.630000 ;
      RECT 873.790000 0.000000 877.875000 0.630000 ;
      RECT 869.290000 0.000000 873.370000 0.630000 ;
      RECT 864.785000 0.000000 868.870000 0.630000 ;
      RECT 860.285000 0.000000 864.365000 0.630000 ;
      RECT 855.780000 0.000000 859.865000 0.630000 ;
      RECT 851.275000 0.000000 855.360000 0.630000 ;
      RECT 846.775000 0.000000 850.855000 0.630000 ;
      RECT 842.270000 0.000000 846.355000 0.630000 ;
      RECT 837.770000 0.000000 841.850000 0.630000 ;
      RECT 833.265000 0.000000 837.350000 0.630000 ;
      RECT 828.760000 0.000000 832.845000 0.630000 ;
      RECT 824.260000 0.000000 828.340000 0.630000 ;
      RECT 819.755000 0.000000 823.840000 0.630000 ;
      RECT 815.255000 0.000000 819.335000 0.630000 ;
      RECT 810.750000 0.000000 814.835000 0.630000 ;
      RECT 806.245000 0.000000 810.330000 0.630000 ;
      RECT 801.745000 0.000000 805.825000 0.630000 ;
      RECT 797.240000 0.000000 801.325000 0.630000 ;
      RECT 792.740000 0.000000 796.820000 0.630000 ;
      RECT 788.235000 0.000000 792.320000 0.630000 ;
      RECT 783.730000 0.000000 787.815000 0.630000 ;
      RECT 779.230000 0.000000 783.310000 0.630000 ;
      RECT 774.725000 0.000000 778.810000 0.630000 ;
      RECT 770.225000 0.000000 774.305000 0.630000 ;
      RECT 765.720000 0.000000 769.805000 0.630000 ;
      RECT 761.215000 0.000000 765.300000 0.630000 ;
      RECT 756.715000 0.000000 760.795000 0.630000 ;
      RECT 752.210000 0.000000 756.295000 0.630000 ;
      RECT 747.710000 0.000000 751.790000 0.630000 ;
      RECT 743.205000 0.000000 747.290000 0.630000 ;
      RECT 738.700000 0.000000 742.785000 0.630000 ;
      RECT 734.200000 0.000000 738.280000 0.630000 ;
      RECT 729.695000 0.000000 733.780000 0.630000 ;
      RECT 725.195000 0.000000 729.275000 0.630000 ;
      RECT 720.690000 0.000000 724.775000 0.630000 ;
      RECT 716.185000 0.000000 720.270000 0.630000 ;
      RECT 711.685000 0.000000 715.765000 0.630000 ;
      RECT 707.180000 0.000000 711.265000 0.630000 ;
      RECT 702.680000 0.000000 706.760000 0.630000 ;
      RECT 698.175000 0.000000 702.260000 0.630000 ;
      RECT 693.670000 0.000000 697.755000 0.630000 ;
      RECT 689.170000 0.000000 693.250000 0.630000 ;
      RECT 684.665000 0.000000 688.750000 0.630000 ;
      RECT 680.165000 0.000000 684.245000 0.630000 ;
      RECT 675.660000 0.000000 679.745000 0.630000 ;
      RECT 671.155000 0.000000 675.240000 0.630000 ;
      RECT 666.655000 0.000000 670.735000 0.630000 ;
      RECT 662.150000 0.000000 666.235000 0.630000 ;
      RECT 657.650000 0.000000 661.730000 0.630000 ;
      RECT 653.145000 0.000000 657.230000 0.630000 ;
      RECT 648.640000 0.000000 652.725000 0.630000 ;
      RECT 644.140000 0.000000 648.220000 0.630000 ;
      RECT 639.635000 0.000000 643.720000 0.630000 ;
      RECT 635.135000 0.000000 639.215000 0.630000 ;
      RECT 630.630000 0.000000 634.715000 0.630000 ;
      RECT 626.125000 0.000000 630.210000 0.630000 ;
      RECT 621.625000 0.000000 625.705000 0.630000 ;
      RECT 617.120000 0.000000 621.205000 0.630000 ;
      RECT 612.620000 0.000000 616.700000 0.630000 ;
      RECT 608.115000 0.000000 612.200000 0.630000 ;
      RECT 603.610000 0.000000 607.695000 0.630000 ;
      RECT 599.110000 0.000000 603.190000 0.630000 ;
      RECT 594.605000 0.000000 598.690000 0.630000 ;
      RECT 590.105000 0.000000 594.185000 0.630000 ;
      RECT 585.600000 0.000000 589.685000 0.630000 ;
      RECT 581.095000 0.000000 585.180000 0.630000 ;
      RECT 576.595000 0.000000 580.675000 0.630000 ;
      RECT 572.090000 0.000000 576.175000 0.630000 ;
      RECT 567.590000 0.000000 571.670000 0.630000 ;
      RECT 563.085000 0.000000 567.170000 0.630000 ;
      RECT 558.580000 0.000000 562.665000 0.630000 ;
      RECT 554.080000 0.000000 558.160000 0.630000 ;
      RECT 549.575000 0.000000 553.660000 0.630000 ;
      RECT 545.075000 0.000000 549.155000 0.630000 ;
      RECT 540.570000 0.000000 544.655000 0.630000 ;
      RECT 536.065000 0.000000 540.150000 0.630000 ;
      RECT 531.565000 0.000000 535.645000 0.630000 ;
      RECT 527.060000 0.000000 531.145000 0.630000 ;
      RECT 522.560000 0.000000 526.640000 0.630000 ;
      RECT 518.055000 0.000000 522.140000 0.630000 ;
      RECT 513.550000 0.000000 517.635000 0.630000 ;
      RECT 509.050000 0.000000 513.130000 0.630000 ;
      RECT 504.545000 0.000000 508.630000 0.630000 ;
      RECT 500.045000 0.000000 504.125000 0.630000 ;
      RECT 495.540000 0.000000 499.625000 0.630000 ;
      RECT 491.035000 0.000000 495.120000 0.630000 ;
      RECT 486.535000 0.000000 490.615000 0.630000 ;
      RECT 482.030000 0.000000 486.115000 0.630000 ;
      RECT 477.530000 0.000000 481.610000 0.630000 ;
      RECT 473.025000 0.000000 477.110000 0.630000 ;
      RECT 468.520000 0.000000 472.605000 0.630000 ;
      RECT 464.020000 0.000000 468.100000 0.630000 ;
      RECT 459.515000 0.000000 463.600000 0.630000 ;
      RECT 455.015000 0.000000 459.095000 0.630000 ;
      RECT 450.510000 0.000000 454.595000 0.630000 ;
      RECT 446.005000 0.000000 450.090000 0.630000 ;
      RECT 441.505000 0.000000 445.585000 0.630000 ;
      RECT 437.000000 0.000000 441.085000 0.630000 ;
      RECT 432.500000 0.000000 436.580000 0.630000 ;
      RECT 427.995000 0.000000 432.080000 0.630000 ;
      RECT 423.490000 0.000000 427.575000 0.630000 ;
      RECT 418.990000 0.000000 423.070000 0.630000 ;
      RECT 414.485000 0.000000 418.570000 0.630000 ;
      RECT 409.985000 0.000000 414.065000 0.630000 ;
      RECT 405.480000 0.000000 409.565000 0.630000 ;
      RECT 400.975000 0.000000 405.060000 0.630000 ;
      RECT 396.475000 0.000000 400.555000 0.630000 ;
      RECT 391.970000 0.000000 396.055000 0.630000 ;
      RECT 387.470000 0.000000 391.550000 0.630000 ;
      RECT 382.965000 0.000000 387.050000 0.630000 ;
      RECT 378.460000 0.000000 382.545000 0.630000 ;
      RECT 373.960000 0.000000 378.040000 0.630000 ;
      RECT 369.455000 0.000000 373.540000 0.630000 ;
      RECT 364.955000 0.000000 369.035000 0.630000 ;
      RECT 360.450000 0.000000 364.535000 0.630000 ;
      RECT 355.945000 0.000000 360.030000 0.630000 ;
      RECT 351.445000 0.000000 355.525000 0.630000 ;
      RECT 346.940000 0.000000 351.025000 0.630000 ;
      RECT 342.440000 0.000000 346.520000 0.630000 ;
      RECT 337.935000 0.000000 342.020000 0.630000 ;
      RECT 333.430000 0.000000 337.515000 0.630000 ;
      RECT 328.930000 0.000000 333.010000 0.630000 ;
      RECT 324.425000 0.000000 328.510000 0.630000 ;
      RECT 319.925000 0.000000 324.005000 0.630000 ;
      RECT 315.420000 0.000000 319.505000 0.630000 ;
      RECT 310.915000 0.000000 315.000000 0.630000 ;
      RECT 306.415000 0.000000 310.495000 0.630000 ;
      RECT 301.910000 0.000000 305.995000 0.630000 ;
      RECT 297.410000 0.000000 301.490000 0.630000 ;
      RECT 292.905000 0.000000 296.990000 0.630000 ;
      RECT 288.400000 0.000000 292.485000 0.630000 ;
      RECT 283.900000 0.000000 287.980000 0.630000 ;
      RECT 279.395000 0.000000 283.480000 0.630000 ;
      RECT 274.895000 0.000000 278.975000 0.630000 ;
      RECT 270.390000 0.000000 274.475000 0.630000 ;
      RECT 265.885000 0.000000 269.970000 0.630000 ;
      RECT 261.385000 0.000000 265.465000 0.630000 ;
      RECT 256.880000 0.000000 260.965000 0.630000 ;
      RECT 252.380000 0.000000 256.460000 0.630000 ;
      RECT 247.875000 0.000000 251.960000 0.630000 ;
      RECT 243.370000 0.000000 247.455000 0.630000 ;
      RECT 238.870000 0.000000 242.950000 0.630000 ;
      RECT 234.365000 0.000000 238.450000 0.630000 ;
      RECT 229.865000 0.000000 233.945000 0.630000 ;
      RECT 225.360000 0.000000 229.445000 0.630000 ;
      RECT 220.855000 0.000000 224.940000 0.630000 ;
      RECT 216.355000 0.000000 220.435000 0.630000 ;
      RECT 211.850000 0.000000 215.935000 0.630000 ;
      RECT 207.350000 0.000000 211.430000 0.630000 ;
      RECT 202.845000 0.000000 206.930000 0.630000 ;
      RECT 198.340000 0.000000 202.425000 0.630000 ;
      RECT 193.840000 0.000000 197.920000 0.630000 ;
      RECT 189.335000 0.000000 193.420000 0.630000 ;
      RECT 184.835000 0.000000 188.915000 0.630000 ;
      RECT 180.330000 0.000000 184.415000 0.630000 ;
      RECT 175.825000 0.000000 179.910000 0.630000 ;
      RECT 171.325000 0.000000 175.405000 0.630000 ;
      RECT 166.820000 0.000000 170.905000 0.630000 ;
      RECT 162.320000 0.000000 166.400000 0.630000 ;
      RECT 157.815000 0.000000 161.900000 0.630000 ;
      RECT 153.310000 0.000000 157.395000 0.630000 ;
      RECT 148.810000 0.000000 152.890000 0.630000 ;
      RECT 144.305000 0.000000 148.390000 0.630000 ;
      RECT 139.805000 0.000000 143.885000 0.630000 ;
      RECT 135.300000 0.000000 139.385000 0.630000 ;
      RECT 130.795000 0.000000 134.880000 0.630000 ;
      RECT 126.295000 0.000000 130.375000 0.630000 ;
      RECT 121.790000 0.000000 125.875000 0.630000 ;
      RECT 117.290000 0.000000 121.370000 0.630000 ;
      RECT 112.785000 0.000000 116.870000 0.630000 ;
      RECT 108.280000 0.000000 112.365000 0.630000 ;
      RECT 103.780000 0.000000 107.860000 0.630000 ;
      RECT 99.275000 0.000000 103.360000 0.630000 ;
      RECT 94.775000 0.000000 98.855000 0.630000 ;
      RECT 90.270000 0.000000 94.355000 0.630000 ;
      RECT 85.765000 0.000000 89.850000 0.630000 ;
      RECT 81.265000 0.000000 85.345000 0.630000 ;
      RECT 76.760000 0.000000 80.845000 0.630000 ;
      RECT 72.260000 0.000000 76.340000 0.630000 ;
      RECT 67.755000 0.000000 71.840000 0.630000 ;
      RECT 63.250000 0.000000 67.335000 0.630000 ;
      RECT 58.750000 0.000000 62.830000 0.630000 ;
      RECT 54.245000 0.000000 58.330000 0.630000 ;
      RECT 49.745000 0.000000 53.825000 0.630000 ;
      RECT 45.240000 0.000000 49.325000 0.630000 ;
      RECT 40.735000 0.000000 44.820000 0.630000 ;
      RECT 36.235000 0.000000 40.315000 0.630000 ;
      RECT 31.730000 0.000000 35.815000 0.630000 ;
      RECT 27.230000 0.000000 31.310000 0.630000 ;
      RECT 22.725000 0.000000 26.810000 0.630000 ;
      RECT 18.220000 0.000000 22.305000 0.630000 ;
      RECT 13.720000 0.000000 17.800000 0.630000 ;
      RECT 9.215000 0.000000 13.300000 0.630000 ;
      RECT 4.715000 0.000000 8.795000 0.630000 ;
      RECT 1.820000 0.000000 4.295000 0.630000 ;
      RECT 0.000000 0.000000 1.400000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 2936.040000 2220.420000 2939.640000 ;
      RECT 1.100000 2935.430000 2220.420000 2936.040000 ;
      RECT 1.100000 2935.140000 2219.320000 2935.430000 ;
      RECT 0.000000 2934.530000 2219.320000 2935.140000 ;
      RECT 0.000000 2884.580000 2220.420000 2934.530000 ;
      RECT 1.100000 2883.680000 2220.420000 2884.580000 ;
      RECT 0.000000 2883.530000 2220.420000 2883.680000 ;
      RECT 0.000000 2882.630000 2219.320000 2883.530000 ;
      RECT 0.000000 2829.115000 2220.420000 2882.630000 ;
      RECT 1.100000 2828.215000 2220.420000 2829.115000 ;
      RECT 0.000000 2827.000000 2220.420000 2828.215000 ;
      RECT 0.000000 2826.100000 2219.320000 2827.000000 ;
      RECT 0.000000 2773.650000 2220.420000 2826.100000 ;
      RECT 1.100000 2772.750000 2220.420000 2773.650000 ;
      RECT 0.000000 2770.470000 2220.420000 2772.750000 ;
      RECT 0.000000 2769.570000 2219.320000 2770.470000 ;
      RECT 0.000000 2718.185000 2220.420000 2769.570000 ;
      RECT 1.100000 2717.285000 2220.420000 2718.185000 ;
      RECT 0.000000 2713.940000 2220.420000 2717.285000 ;
      RECT 0.000000 2713.040000 2219.320000 2713.940000 ;
      RECT 0.000000 2662.720000 2220.420000 2713.040000 ;
      RECT 1.100000 2661.820000 2220.420000 2662.720000 ;
      RECT 0.000000 2657.405000 2220.420000 2661.820000 ;
      RECT 0.000000 2656.505000 2219.320000 2657.405000 ;
      RECT 0.000000 2607.260000 2220.420000 2656.505000 ;
      RECT 1.100000 2606.360000 2220.420000 2607.260000 ;
      RECT 0.000000 2600.875000 2220.420000 2606.360000 ;
      RECT 0.000000 2599.975000 2219.320000 2600.875000 ;
      RECT 0.000000 2551.795000 2220.420000 2599.975000 ;
      RECT 1.100000 2550.895000 2220.420000 2551.795000 ;
      RECT 0.000000 2544.345000 2220.420000 2550.895000 ;
      RECT 0.000000 2543.445000 2219.320000 2544.345000 ;
      RECT 0.000000 2496.330000 2220.420000 2543.445000 ;
      RECT 1.100000 2495.430000 2220.420000 2496.330000 ;
      RECT 0.000000 2487.815000 2220.420000 2495.430000 ;
      RECT 0.000000 2486.915000 2219.320000 2487.815000 ;
      RECT 0.000000 2440.865000 2220.420000 2486.915000 ;
      RECT 1.100000 2439.965000 2220.420000 2440.865000 ;
      RECT 0.000000 2431.285000 2220.420000 2439.965000 ;
      RECT 0.000000 2430.385000 2219.320000 2431.285000 ;
      RECT 0.000000 2385.400000 2220.420000 2430.385000 ;
      RECT 1.100000 2384.500000 2220.420000 2385.400000 ;
      RECT 0.000000 2374.750000 2220.420000 2384.500000 ;
      RECT 0.000000 2373.850000 2219.320000 2374.750000 ;
      RECT 0.000000 2329.940000 2220.420000 2373.850000 ;
      RECT 1.100000 2329.040000 2220.420000 2329.940000 ;
      RECT 0.000000 2318.220000 2220.420000 2329.040000 ;
      RECT 0.000000 2317.320000 2219.320000 2318.220000 ;
      RECT 0.000000 2274.475000 2220.420000 2317.320000 ;
      RECT 1.100000 2273.575000 2220.420000 2274.475000 ;
      RECT 0.000000 2261.690000 2220.420000 2273.575000 ;
      RECT 0.000000 2260.790000 2219.320000 2261.690000 ;
      RECT 0.000000 2219.010000 2220.420000 2260.790000 ;
      RECT 1.100000 2218.110000 2220.420000 2219.010000 ;
      RECT 0.000000 2205.160000 2220.420000 2218.110000 ;
      RECT 0.000000 2204.260000 2219.320000 2205.160000 ;
      RECT 0.000000 2163.545000 2220.420000 2204.260000 ;
      RECT 1.100000 2162.645000 2220.420000 2163.545000 ;
      RECT 0.000000 2148.630000 2220.420000 2162.645000 ;
      RECT 0.000000 2147.730000 2219.320000 2148.630000 ;
      RECT 0.000000 2108.080000 2220.420000 2147.730000 ;
      RECT 1.100000 2107.180000 2220.420000 2108.080000 ;
      RECT 0.000000 2092.095000 2220.420000 2107.180000 ;
      RECT 0.000000 2091.195000 2219.320000 2092.095000 ;
      RECT 0.000000 2052.620000 2220.420000 2091.195000 ;
      RECT 1.100000 2051.720000 2220.420000 2052.620000 ;
      RECT 0.000000 2035.565000 2220.420000 2051.720000 ;
      RECT 0.000000 2034.665000 2219.320000 2035.565000 ;
      RECT 0.000000 1997.155000 2220.420000 2034.665000 ;
      RECT 1.100000 1996.255000 2220.420000 1997.155000 ;
      RECT 0.000000 1979.035000 2220.420000 1996.255000 ;
      RECT 0.000000 1978.135000 2219.320000 1979.035000 ;
      RECT 0.000000 1941.690000 2220.420000 1978.135000 ;
      RECT 1.100000 1940.790000 2220.420000 1941.690000 ;
      RECT 0.000000 1922.505000 2220.420000 1940.790000 ;
      RECT 0.000000 1921.605000 2219.320000 1922.505000 ;
      RECT 0.000000 1886.225000 2220.420000 1921.605000 ;
      RECT 1.100000 1885.325000 2220.420000 1886.225000 ;
      RECT 0.000000 1865.975000 2220.420000 1885.325000 ;
      RECT 0.000000 1865.075000 2219.320000 1865.975000 ;
      RECT 0.000000 1830.760000 2220.420000 1865.075000 ;
      RECT 1.100000 1829.860000 2220.420000 1830.760000 ;
      RECT 0.000000 1809.440000 2220.420000 1829.860000 ;
      RECT 0.000000 1808.540000 2219.320000 1809.440000 ;
      RECT 0.000000 1775.300000 2220.420000 1808.540000 ;
      RECT 1.100000 1774.400000 2220.420000 1775.300000 ;
      RECT 0.000000 1752.910000 2220.420000 1774.400000 ;
      RECT 0.000000 1752.010000 2219.320000 1752.910000 ;
      RECT 0.000000 1719.835000 2220.420000 1752.010000 ;
      RECT 1.100000 1718.935000 2220.420000 1719.835000 ;
      RECT 0.000000 1696.380000 2220.420000 1718.935000 ;
      RECT 0.000000 1695.480000 2219.320000 1696.380000 ;
      RECT 0.000000 1664.370000 2220.420000 1695.480000 ;
      RECT 1.100000 1663.470000 2220.420000 1664.370000 ;
      RECT 0.000000 1639.850000 2220.420000 1663.470000 ;
      RECT 0.000000 1638.950000 2219.320000 1639.850000 ;
      RECT 0.000000 1608.905000 2220.420000 1638.950000 ;
      RECT 1.100000 1608.005000 2220.420000 1608.905000 ;
      RECT 0.000000 1583.320000 2220.420000 1608.005000 ;
      RECT 0.000000 1582.420000 2219.320000 1583.320000 ;
      RECT 0.000000 1553.440000 2220.420000 1582.420000 ;
      RECT 1.100000 1552.540000 2220.420000 1553.440000 ;
      RECT 0.000000 1526.785000 2220.420000 1552.540000 ;
      RECT 0.000000 1525.885000 2219.320000 1526.785000 ;
      RECT 0.000000 1497.980000 2220.420000 1525.885000 ;
      RECT 1.100000 1497.080000 2220.420000 1497.980000 ;
      RECT 0.000000 1470.255000 2220.420000 1497.080000 ;
      RECT 0.000000 1469.355000 2219.320000 1470.255000 ;
      RECT 0.000000 1442.515000 2220.420000 1469.355000 ;
      RECT 1.100000 1441.615000 2220.420000 1442.515000 ;
      RECT 0.000000 1413.725000 2220.420000 1441.615000 ;
      RECT 0.000000 1412.825000 2219.320000 1413.725000 ;
      RECT 0.000000 1387.050000 2220.420000 1412.825000 ;
      RECT 1.100000 1386.150000 2220.420000 1387.050000 ;
      RECT 0.000000 1357.195000 2220.420000 1386.150000 ;
      RECT 0.000000 1356.295000 2219.320000 1357.195000 ;
      RECT 0.000000 1331.585000 2220.420000 1356.295000 ;
      RECT 1.100000 1330.685000 2220.420000 1331.585000 ;
      RECT 0.000000 1300.665000 2220.420000 1330.685000 ;
      RECT 0.000000 1299.765000 2219.320000 1300.665000 ;
      RECT 0.000000 1276.120000 2220.420000 1299.765000 ;
      RECT 1.100000 1275.220000 2220.420000 1276.120000 ;
      RECT 0.000000 1244.130000 2220.420000 1275.220000 ;
      RECT 0.000000 1243.230000 2219.320000 1244.130000 ;
      RECT 0.000000 1220.660000 2220.420000 1243.230000 ;
      RECT 1.100000 1219.760000 2220.420000 1220.660000 ;
      RECT 0.000000 1187.600000 2220.420000 1219.760000 ;
      RECT 0.000000 1186.700000 2219.320000 1187.600000 ;
      RECT 0.000000 1165.195000 2220.420000 1186.700000 ;
      RECT 1.100000 1164.295000 2220.420000 1165.195000 ;
      RECT 0.000000 1131.070000 2220.420000 1164.295000 ;
      RECT 0.000000 1130.170000 2219.320000 1131.070000 ;
      RECT 0.000000 1109.730000 2220.420000 1130.170000 ;
      RECT 1.100000 1108.830000 2220.420000 1109.730000 ;
      RECT 0.000000 1074.540000 2220.420000 1108.830000 ;
      RECT 0.000000 1073.640000 2219.320000 1074.540000 ;
      RECT 0.000000 1054.265000 2220.420000 1073.640000 ;
      RECT 1.100000 1053.365000 2220.420000 1054.265000 ;
      RECT 0.000000 1018.010000 2220.420000 1053.365000 ;
      RECT 0.000000 1017.110000 2219.320000 1018.010000 ;
      RECT 0.000000 998.800000 2220.420000 1017.110000 ;
      RECT 1.100000 997.900000 2220.420000 998.800000 ;
      RECT 0.000000 961.475000 2220.420000 997.900000 ;
      RECT 0.000000 960.575000 2219.320000 961.475000 ;
      RECT 0.000000 943.340000 2220.420000 960.575000 ;
      RECT 1.100000 942.440000 2220.420000 943.340000 ;
      RECT 0.000000 904.945000 2220.420000 942.440000 ;
      RECT 0.000000 904.045000 2219.320000 904.945000 ;
      RECT 0.000000 887.875000 2220.420000 904.045000 ;
      RECT 1.100000 886.975000 2220.420000 887.875000 ;
      RECT 0.000000 848.415000 2220.420000 886.975000 ;
      RECT 0.000000 847.515000 2219.320000 848.415000 ;
      RECT 0.000000 832.410000 2220.420000 847.515000 ;
      RECT 1.100000 831.510000 2220.420000 832.410000 ;
      RECT 0.000000 791.885000 2220.420000 831.510000 ;
      RECT 0.000000 790.985000 2219.320000 791.885000 ;
      RECT 0.000000 776.945000 2220.420000 790.985000 ;
      RECT 1.100000 776.045000 2220.420000 776.945000 ;
      RECT 0.000000 735.355000 2220.420000 776.045000 ;
      RECT 0.000000 734.455000 2219.320000 735.355000 ;
      RECT 0.000000 721.480000 2220.420000 734.455000 ;
      RECT 1.100000 720.580000 2220.420000 721.480000 ;
      RECT 0.000000 678.820000 2220.420000 720.580000 ;
      RECT 0.000000 677.920000 2219.320000 678.820000 ;
      RECT 0.000000 666.020000 2220.420000 677.920000 ;
      RECT 1.100000 665.120000 2220.420000 666.020000 ;
      RECT 0.000000 622.290000 2220.420000 665.120000 ;
      RECT 0.000000 621.390000 2219.320000 622.290000 ;
      RECT 0.000000 610.555000 2220.420000 621.390000 ;
      RECT 1.100000 609.655000 2220.420000 610.555000 ;
      RECT 0.000000 565.760000 2220.420000 609.655000 ;
      RECT 0.000000 564.860000 2219.320000 565.760000 ;
      RECT 0.000000 555.090000 2220.420000 564.860000 ;
      RECT 1.100000 554.190000 2220.420000 555.090000 ;
      RECT 0.000000 509.230000 2220.420000 554.190000 ;
      RECT 0.000000 508.330000 2219.320000 509.230000 ;
      RECT 0.000000 499.625000 2220.420000 508.330000 ;
      RECT 1.100000 498.725000 2220.420000 499.625000 ;
      RECT 0.000000 452.700000 2220.420000 498.725000 ;
      RECT 0.000000 451.800000 2219.320000 452.700000 ;
      RECT 0.000000 444.160000 2220.420000 451.800000 ;
      RECT 1.100000 443.260000 2220.420000 444.160000 ;
      RECT 0.000000 396.165000 2220.420000 443.260000 ;
      RECT 0.000000 395.265000 2219.320000 396.165000 ;
      RECT 0.000000 388.700000 2220.420000 395.265000 ;
      RECT 1.100000 387.800000 2220.420000 388.700000 ;
      RECT 0.000000 339.635000 2220.420000 387.800000 ;
      RECT 0.000000 338.735000 2219.320000 339.635000 ;
      RECT 0.000000 333.235000 2220.420000 338.735000 ;
      RECT 1.100000 332.335000 2220.420000 333.235000 ;
      RECT 0.000000 283.105000 2220.420000 332.335000 ;
      RECT 0.000000 282.205000 2219.320000 283.105000 ;
      RECT 0.000000 277.770000 2220.420000 282.205000 ;
      RECT 1.100000 276.870000 2220.420000 277.770000 ;
      RECT 0.000000 226.575000 2220.420000 276.870000 ;
      RECT 0.000000 225.675000 2219.320000 226.575000 ;
      RECT 0.000000 222.305000 2220.420000 225.675000 ;
      RECT 1.100000 221.405000 2220.420000 222.305000 ;
      RECT 0.000000 170.045000 2220.420000 221.405000 ;
      RECT 0.000000 169.145000 2219.320000 170.045000 ;
      RECT 0.000000 166.840000 2220.420000 169.145000 ;
      RECT 1.100000 165.940000 2220.420000 166.840000 ;
      RECT 0.000000 113.510000 2220.420000 165.940000 ;
      RECT 0.000000 112.610000 2219.320000 113.510000 ;
      RECT 0.000000 111.380000 2220.420000 112.610000 ;
      RECT 1.100000 110.480000 2220.420000 111.380000 ;
      RECT 0.000000 56.980000 2220.420000 110.480000 ;
      RECT 0.000000 56.080000 2219.320000 56.980000 ;
      RECT 0.000000 55.915000 2220.420000 56.080000 ;
      RECT 1.100000 55.015000 2220.420000 55.915000 ;
      RECT 0.000000 3.770000 2220.420000 55.015000 ;
      RECT 1.100000 3.160000 2220.420000 3.770000 ;
      RECT 1.100000 2.870000 2219.320000 3.160000 ;
      RECT 0.000000 2.260000 2219.320000 2.870000 ;
      RECT 0.000000 0.000000 2220.420000 2.260000 ;
    LAYER met4 ;
      RECT 0.000000 2937.330000 2220.420000 2939.640000 ;
      RECT 4.360000 2933.330000 2216.060000 2937.330000 ;
      RECT 2214.660000 5.630000 2216.060000 2933.330000 ;
      RECT 8.360000 5.630000 2212.060000 2933.330000 ;
      RECT 4.360000 5.630000 5.760000 2933.330000 ;
      RECT 2218.660000 1.630000 2220.420000 2937.330000 ;
      RECT 4.360000 1.630000 2216.060000 5.630000 ;
      RECT 0.000000 1.630000 1.760000 2937.330000 ;
      RECT 0.000000 0.000000 2220.420000 1.630000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
